

module div(
    input wire clock,
    input wire reset,

    input wire in_valid,
    input wire [63:0] in_a,
    input wire [63:0] in_b,
    input wire div_signed,

    output wire result_valid,
    output wire [63:0]quotient,
    output wire [63:0]remainder
);
    


endmodule



