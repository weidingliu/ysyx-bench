module IF(
  input         clock,
  input         reset,
  input         io_branch_io_is_branch,
  input         io_branch_io_is_jump,
  input  [63:0] io_branch_io_dnpc,
  output        io_cache_req_addr_req_valid,
  output [63:0] io_cache_req_addr_req_bits_addr,
  output        io_cache_req_rdata_rep_ready,
  input         io_cache_req_rdata_rep_valid,
  input  [63:0] io_cache_req_rdata_rep_bits_rdata,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_PC,
  output [31:0] io_out_bits_Inst,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] temp; // @[IF.scala 22:21]
  wire [63:0] _temp_T_3 = temp + 64'h4; // @[IF.scala 23:136]
  wire [31:0] inst = temp[2] ? io_cache_req_rdata_rep_bits_rdata[63:32] : io_cache_req_rdata_rep_bits_rdata[31:0]; // @[IF.scala 40:17]
  assign io_cache_req_addr_req_valid = io_out_ready; // @[IF.scala 34:37]
  assign io_cache_req_addr_req_bits_addr = temp; // @[IF.scala 33:35]
  assign io_cache_req_rdata_rep_ready = io_out_ready; // @[IF.scala 39:32]
  assign io_out_valid = io_cache_req_rdata_rep_valid; // @[IF.scala 31:22]
  assign io_out_bits_PC = temp; // @[IF.scala 42:18]
  assign io_out_bits_Inst = io_flush ? 32'h0 : inst; // @[IF.scala 43:26]
  always @(posedge clock) begin
    if (reset) begin // @[IF.scala 22:21]
      temp <= 64'h80000000; // @[IF.scala 22:21]
    end else if (io_branch_io_is_jump | io_branch_io_is_branch) begin // @[IF.scala 23:14]
      temp <= io_branch_io_dnpc;
    end else if (io_out_ready & io_cache_req_rdata_rep_valid) begin // @[IF.scala 23:85]
      temp <= _temp_T_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  temp = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ID(
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_PC,
  input  [31:0] io_in_bits_Inst,
  input  [63:0] io_REG1,
  input  [63:0] io_REG2,
  input         io_flush,
  input         io_out_ready,
  output        io_out_valid,
  output [2:0]  io_out_bits_ctrl_signal_src1Type,
  output [2:0]  io_out_bits_ctrl_signal_src2Type,
  output [2:0]  io_out_bits_ctrl_signal_fuType,
  output        io_out_bits_ctrl_signal_inst_valid,
  output [4:0]  io_out_bits_ctrl_signal_rfSrc1,
  output [4:0]  io_out_bits_ctrl_signal_rfSrc2,
  output        io_out_bits_ctrl_signal_rfWen,
  output [6:0]  io_out_bits_ctrl_signal_aluoptype,
  output [4:0]  io_out_bits_ctrl_signal_rfDest,
  output [63:0] io_out_bits_ctrl_data_src1,
  output [63:0] io_out_bits_ctrl_data_src2,
  output [63:0] io_out_bits_ctrl_data_Imm,
  output [63:0] io_out_bits_ctrl_flow_PC,
  output [31:0] io_out_bits_ctrl_flow_inst
);
  wire [4:0] rd = io_in_bits_Inst[11:7]; // @[ID.scala 51:88]
  wire [31:0] _Inst_decode_T = io_in_bits_Inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_1 = 32'h13 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire [31:0] _Inst_decode_T_2 = io_in_bits_Inst & 32'hfc00707f; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_3 = 32'h1013 == _Inst_decode_T_2; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_5 = 32'h6013 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_7 = 32'h3003 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_9 = 32'h2003 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_11 = 32'h3013 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_13 = 32'h1b == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_15 = 32'h40005013 == _Inst_decode_T_2; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_17 = 32'h4003 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_19 = 32'h3 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_21 = 32'h4013 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_23 = 32'h7013 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_25 = 32'h5013 == _Inst_decode_T_2; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_27 = 32'h1003 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_29 = 32'h5003 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_31 = 32'h101b == _Inst_decode_T_2; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_33 = 32'h4000501b == _Inst_decode_T_2; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_35 = 32'h501b == _Inst_decode_T_2; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_37 = 32'h2013 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_39 = 32'h6003 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire [31:0] _Inst_decode_T_40 = io_in_bits_Inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_41 = 32'h3b == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_43 = 32'h40000033 == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_45 = 32'h33 == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_47 = 32'h7033 == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_49 = 32'h3033 == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_51 = 32'h103b == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_53 = 32'h6033 == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_55 = 32'h200003b == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_57 = 32'h200403b == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_59 = 32'h200603b == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_61 = 32'h4000003b == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_63 = 32'h2033 == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_65 = 32'h4000503b == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_67 = 32'h503b == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_69 = 32'h4033 == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_71 = 32'h200703b == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_73 = 32'h1033 == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_75 = 32'h2007033 == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_77 = 32'h200503b == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_79 = 32'h2006033 == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_81 = 32'h5033 == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_83 = 32'h2005033 == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_85 = 32'h2004033 == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_87 = 32'h40005033 == _Inst_decode_T_2; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_89 = 32'h2000033 == _Inst_decode_T_40; // @[Lookup.scala 31:38]
  wire [31:0] _Inst_decode_T_90 = io_in_bits_Inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_91 = 32'h17 == _Inst_decode_T_90; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_93 = 32'h37 == _Inst_decode_T_90; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_95 = 32'h3023 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_97 = 32'h1023 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_99 = 32'h23 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_101 = 32'h2023 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_103 = 32'h100073 == io_in_bits_Inst; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_105 = 32'h6f == _Inst_decode_T_90; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_107 = 32'h67 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_109 = 32'h63 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_111 = 32'h1063 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_113 = 32'h5063 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_115 = 32'h4063 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_117 = 32'h6063 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_119 = 32'h7063 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_121 = 32'h2073 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_123 = 32'h1073 == _Inst_decode_T; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_125 = 32'h73 == io_in_bits_Inst; // @[Lookup.scala 31:38]
  wire  _Inst_decode_T_127 = 32'h30200073 == io_in_bits_Inst; // @[Lookup.scala 31:38]
  wire [3:0] _Inst_decode_T_130 = _Inst_decode_T_123 ? 4'h8 : 4'h0; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_131 = _Inst_decode_T_121 ? 4'h8 : _Inst_decode_T_130; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_132 = _Inst_decode_T_119 ? 4'hb : _Inst_decode_T_131; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_133 = _Inst_decode_T_117 ? 4'hb : _Inst_decode_T_132; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_134 = _Inst_decode_T_115 ? 4'hb : _Inst_decode_T_133; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_135 = _Inst_decode_T_113 ? 4'hb : _Inst_decode_T_134; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_136 = _Inst_decode_T_111 ? 4'hb : _Inst_decode_T_135; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_137 = _Inst_decode_T_109 ? 4'hb : _Inst_decode_T_136; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_138 = _Inst_decode_T_107 ? 4'h8 : _Inst_decode_T_137; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_139 = _Inst_decode_T_105 ? 4'h7 : _Inst_decode_T_138; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_140 = _Inst_decode_T_103 ? 4'h0 : _Inst_decode_T_139; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_141 = _Inst_decode_T_101 ? 4'h9 : _Inst_decode_T_140; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_142 = _Inst_decode_T_99 ? 4'h9 : _Inst_decode_T_141; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_143 = _Inst_decode_T_97 ? 4'h9 : _Inst_decode_T_142; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_144 = _Inst_decode_T_95 ? 4'h9 : _Inst_decode_T_143; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_145 = _Inst_decode_T_93 ? 4'h3 : _Inst_decode_T_144; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_146 = _Inst_decode_T_91 ? 4'h3 : _Inst_decode_T_145; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_147 = _Inst_decode_T_89 ? 4'h5 : _Inst_decode_T_146; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_148 = _Inst_decode_T_87 ? 4'h5 : _Inst_decode_T_147; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_149 = _Inst_decode_T_85 ? 4'h5 : _Inst_decode_T_148; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_150 = _Inst_decode_T_83 ? 4'h5 : _Inst_decode_T_149; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_151 = _Inst_decode_T_81 ? 4'h5 : _Inst_decode_T_150; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_152 = _Inst_decode_T_79 ? 4'h5 : _Inst_decode_T_151; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_153 = _Inst_decode_T_77 ? 4'h5 : _Inst_decode_T_152; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_154 = _Inst_decode_T_75 ? 4'h5 : _Inst_decode_T_153; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_155 = _Inst_decode_T_73 ? 4'h5 : _Inst_decode_T_154; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_156 = _Inst_decode_T_71 ? 4'h5 : _Inst_decode_T_155; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_157 = _Inst_decode_T_69 ? 4'h5 : _Inst_decode_T_156; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_158 = _Inst_decode_T_67 ? 4'h5 : _Inst_decode_T_157; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_159 = _Inst_decode_T_65 ? 4'h5 : _Inst_decode_T_158; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_160 = _Inst_decode_T_63 ? 4'h5 : _Inst_decode_T_159; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_161 = _Inst_decode_T_61 ? 4'h5 : _Inst_decode_T_160; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_162 = _Inst_decode_T_59 ? 4'h5 : _Inst_decode_T_161; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_163 = _Inst_decode_T_57 ? 4'h5 : _Inst_decode_T_162; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_164 = _Inst_decode_T_55 ? 4'h5 : _Inst_decode_T_163; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_165 = _Inst_decode_T_53 ? 4'h5 : _Inst_decode_T_164; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_166 = _Inst_decode_T_51 ? 4'h5 : _Inst_decode_T_165; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_167 = _Inst_decode_T_49 ? 4'h5 : _Inst_decode_T_166; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_168 = _Inst_decode_T_47 ? 4'h5 : _Inst_decode_T_167; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_169 = _Inst_decode_T_45 ? 4'h5 : _Inst_decode_T_168; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_170 = _Inst_decode_T_43 ? 4'h5 : _Inst_decode_T_169; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_171 = _Inst_decode_T_41 ? 4'h5 : _Inst_decode_T_170; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_172 = _Inst_decode_T_39 ? 4'h8 : _Inst_decode_T_171; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_173 = _Inst_decode_T_37 ? 4'h8 : _Inst_decode_T_172; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_174 = _Inst_decode_T_35 ? 4'h8 : _Inst_decode_T_173; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_175 = _Inst_decode_T_33 ? 4'h8 : _Inst_decode_T_174; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_176 = _Inst_decode_T_31 ? 4'h8 : _Inst_decode_T_175; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_177 = _Inst_decode_T_29 ? 4'h8 : _Inst_decode_T_176; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_178 = _Inst_decode_T_27 ? 4'h8 : _Inst_decode_T_177; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_179 = _Inst_decode_T_25 ? 4'h8 : _Inst_decode_T_178; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_180 = _Inst_decode_T_23 ? 4'h8 : _Inst_decode_T_179; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_181 = _Inst_decode_T_21 ? 4'h8 : _Inst_decode_T_180; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_182 = _Inst_decode_T_19 ? 4'h8 : _Inst_decode_T_181; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_183 = _Inst_decode_T_17 ? 4'h8 : _Inst_decode_T_182; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_184 = _Inst_decode_T_15 ? 4'h8 : _Inst_decode_T_183; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_185 = _Inst_decode_T_13 ? 4'h8 : _Inst_decode_T_184; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_186 = _Inst_decode_T_11 ? 4'h8 : _Inst_decode_T_185; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_187 = _Inst_decode_T_9 ? 4'h8 : _Inst_decode_T_186; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_188 = _Inst_decode_T_7 ? 4'h8 : _Inst_decode_T_187; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_189 = _Inst_decode_T_5 ? 4'h8 : _Inst_decode_T_188; // @[Lookup.scala 34:39]
  wire [3:0] _Inst_decode_T_190 = _Inst_decode_T_3 ? 4'h8 : _Inst_decode_T_189; // @[Lookup.scala 34:39]
  wire [3:0] Inst_decode_0 = _Inst_decode_T_1 ? 4'h8 : _Inst_decode_T_190; // @[Lookup.scala 34:39]
  wire [1:0] _Inst_decode_T_195 = _Inst_decode_T_119 ? 2'h2 : 2'h0; // @[Lookup.scala 34:39]
  wire [1:0] _Inst_decode_T_196 = _Inst_decode_T_117 ? 2'h2 : _Inst_decode_T_195; // @[Lookup.scala 34:39]
  wire [1:0] _Inst_decode_T_197 = _Inst_decode_T_115 ? 2'h2 : _Inst_decode_T_196; // @[Lookup.scala 34:39]
  wire [1:0] _Inst_decode_T_198 = _Inst_decode_T_113 ? 2'h2 : _Inst_decode_T_197; // @[Lookup.scala 34:39]
  wire [1:0] _Inst_decode_T_199 = _Inst_decode_T_111 ? 2'h2 : _Inst_decode_T_198; // @[Lookup.scala 34:39]
  wire [1:0] _Inst_decode_T_200 = _Inst_decode_T_109 ? 2'h2 : _Inst_decode_T_199; // @[Lookup.scala 34:39]
  wire [1:0] _Inst_decode_T_201 = _Inst_decode_T_107 ? 2'h3 : _Inst_decode_T_200; // @[Lookup.scala 34:39]
  wire [1:0] _Inst_decode_T_202 = _Inst_decode_T_105 ? 2'h3 : _Inst_decode_T_201; // @[Lookup.scala 34:39]
  wire [1:0] _Inst_decode_T_203 = _Inst_decode_T_103 ? 2'h0 : _Inst_decode_T_202; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_204 = _Inst_decode_T_101 ? 3'h4 : {{1'd0}, _Inst_decode_T_203}; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_205 = _Inst_decode_T_99 ? 3'h4 : _Inst_decode_T_204; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_206 = _Inst_decode_T_97 ? 3'h4 : _Inst_decode_T_205; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_207 = _Inst_decode_T_95 ? 3'h4 : _Inst_decode_T_206; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_208 = _Inst_decode_T_93 ? 3'h0 : _Inst_decode_T_207; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_209 = _Inst_decode_T_91 ? 3'h0 : _Inst_decode_T_208; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_210 = _Inst_decode_T_89 ? 3'h0 : _Inst_decode_T_209; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_211 = _Inst_decode_T_87 ? 3'h0 : _Inst_decode_T_210; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_212 = _Inst_decode_T_85 ? 3'h0 : _Inst_decode_T_211; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_213 = _Inst_decode_T_83 ? 3'h0 : _Inst_decode_T_212; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_214 = _Inst_decode_T_81 ? 3'h1 : _Inst_decode_T_213; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_215 = _Inst_decode_T_79 ? 3'h0 : _Inst_decode_T_214; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_216 = _Inst_decode_T_77 ? 3'h0 : _Inst_decode_T_215; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_217 = _Inst_decode_T_75 ? 3'h0 : _Inst_decode_T_216; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_218 = _Inst_decode_T_73 ? 3'h1 : _Inst_decode_T_217; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_219 = _Inst_decode_T_71 ? 3'h0 : _Inst_decode_T_218; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_220 = _Inst_decode_T_69 ? 3'h0 : _Inst_decode_T_219; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_221 = _Inst_decode_T_67 ? 3'h1 : _Inst_decode_T_220; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_222 = _Inst_decode_T_65 ? 3'h1 : _Inst_decode_T_221; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_223 = _Inst_decode_T_63 ? 3'h5 : _Inst_decode_T_222; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_224 = _Inst_decode_T_61 ? 3'h0 : _Inst_decode_T_223; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_225 = _Inst_decode_T_59 ? 3'h0 : _Inst_decode_T_224; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_226 = _Inst_decode_T_57 ? 3'h0 : _Inst_decode_T_225; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_227 = _Inst_decode_T_55 ? 3'h0 : _Inst_decode_T_226; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_228 = _Inst_decode_T_53 ? 3'h0 : _Inst_decode_T_227; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_229 = _Inst_decode_T_51 ? 3'h1 : _Inst_decode_T_228; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_230 = _Inst_decode_T_49 ? 3'h5 : _Inst_decode_T_229; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_231 = _Inst_decode_T_47 ? 3'h0 : _Inst_decode_T_230; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_232 = _Inst_decode_T_45 ? 3'h0 : _Inst_decode_T_231; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_233 = _Inst_decode_T_43 ? 3'h0 : _Inst_decode_T_232; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_234 = _Inst_decode_T_41 ? 3'h0 : _Inst_decode_T_233; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_235 = _Inst_decode_T_39 ? 3'h4 : _Inst_decode_T_234; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_236 = _Inst_decode_T_37 ? 3'h5 : _Inst_decode_T_235; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_237 = _Inst_decode_T_35 ? 3'h1 : _Inst_decode_T_236; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_238 = _Inst_decode_T_33 ? 3'h1 : _Inst_decode_T_237; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_239 = _Inst_decode_T_31 ? 3'h1 : _Inst_decode_T_238; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_240 = _Inst_decode_T_29 ? 3'h4 : _Inst_decode_T_239; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_241 = _Inst_decode_T_27 ? 3'h4 : _Inst_decode_T_240; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_242 = _Inst_decode_T_25 ? 3'h1 : _Inst_decode_T_241; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_243 = _Inst_decode_T_23 ? 3'h0 : _Inst_decode_T_242; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_244 = _Inst_decode_T_21 ? 3'h0 : _Inst_decode_T_243; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_245 = _Inst_decode_T_19 ? 3'h4 : _Inst_decode_T_244; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_246 = _Inst_decode_T_17 ? 3'h4 : _Inst_decode_T_245; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_247 = _Inst_decode_T_15 ? 3'h1 : _Inst_decode_T_246; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_248 = _Inst_decode_T_13 ? 3'h0 : _Inst_decode_T_247; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_249 = _Inst_decode_T_11 ? 3'h5 : _Inst_decode_T_248; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_250 = _Inst_decode_T_9 ? 3'h4 : _Inst_decode_T_249; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_251 = _Inst_decode_T_7 ? 3'h4 : _Inst_decode_T_250; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_252 = _Inst_decode_T_5 ? 3'h0 : _Inst_decode_T_251; // @[Lookup.scala 34:39]
  wire [2:0] _Inst_decode_T_253 = _Inst_decode_T_3 ? 3'h1 : _Inst_decode_T_252; // @[Lookup.scala 34:39]
  wire [4:0] _Inst_decode_T_254 = _Inst_decode_T_127 ? 5'h18 : 5'h0; // @[Lookup.scala 34:39]
  wire [4:0] _Inst_decode_T_255 = _Inst_decode_T_125 ? 5'h17 : _Inst_decode_T_254; // @[Lookup.scala 34:39]
  wire [4:0] _Inst_decode_T_256 = _Inst_decode_T_123 ? 5'h16 : _Inst_decode_T_255; // @[Lookup.scala 34:39]
  wire [4:0] _Inst_decode_T_257 = _Inst_decode_T_121 ? 5'h15 : _Inst_decode_T_256; // @[Lookup.scala 34:39]
  wire [4:0] _Inst_decode_T_258 = _Inst_decode_T_119 ? 5'hc : _Inst_decode_T_257; // @[Lookup.scala 34:39]
  wire [4:0] _Inst_decode_T_259 = _Inst_decode_T_117 ? 5'hb : _Inst_decode_T_258; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_260 = _Inst_decode_T_115 ? 7'h7b : {{2'd0}, _Inst_decode_T_259}; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_261 = _Inst_decode_T_113 ? 7'h76 : _Inst_decode_T_260; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_262 = _Inst_decode_T_111 ? 7'h6c : _Inst_decode_T_261; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_263 = _Inst_decode_T_109 ? 7'h6b : _Inst_decode_T_262; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_264 = _Inst_decode_T_107 ? 7'h48 : _Inst_decode_T_263; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_265 = _Inst_decode_T_105 ? 7'h19 : _Inst_decode_T_264; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_266 = _Inst_decode_T_103 ? 7'h42 : _Inst_decode_T_265; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_267 = _Inst_decode_T_101 ? 7'h77 : _Inst_decode_T_266; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_268 = _Inst_decode_T_99 ? 7'h74 : _Inst_decode_T_267; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_269 = _Inst_decode_T_97 ? 7'h70 : _Inst_decode_T_268; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_270 = _Inst_decode_T_95 ? 7'h46 : _Inst_decode_T_269; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_271 = _Inst_decode_T_93 ? 7'h1a : _Inst_decode_T_270; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_272 = _Inst_decode_T_91 ? 7'h40 : _Inst_decode_T_271; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_273 = _Inst_decode_T_89 ? 7'h7 : _Inst_decode_T_272; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_274 = _Inst_decode_T_87 ? 7'h14 : _Inst_decode_T_273; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_275 = _Inst_decode_T_85 ? 7'h43 : _Inst_decode_T_274; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_276 = _Inst_decode_T_83 ? 7'h13 : _Inst_decode_T_275; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_277 = _Inst_decode_T_81 ? 7'h75 : _Inst_decode_T_276; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_278 = _Inst_decode_T_79 ? 7'h12 : _Inst_decode_T_277; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_279 = _Inst_decode_T_77 ? 7'h10 : _Inst_decode_T_278; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_280 = _Inst_decode_T_75 ? 7'hf : _Inst_decode_T_279; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_281 = _Inst_decode_T_73 ? 7'h41 : _Inst_decode_T_280; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_282 = _Inst_decode_T_71 ? 7'hd : _Inst_decode_T_281; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_283 = _Inst_decode_T_69 ? 7'h72 : _Inst_decode_T_282; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_284 = _Inst_decode_T_67 ? 7'ha : _Inst_decode_T_283; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_285 = _Inst_decode_T_65 ? 7'h9 : _Inst_decode_T_284; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_286 = _Inst_decode_T_63 ? 7'h2 : _Inst_decode_T_285; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_287 = _Inst_decode_T_61 ? 7'h1 : _Inst_decode_T_286; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_288 = _Inst_decode_T_59 ? 7'h7a : _Inst_decode_T_287; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_289 = _Inst_decode_T_57 ? 7'h79 : _Inst_decode_T_288; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_290 = _Inst_decode_T_55 ? 7'h78 : _Inst_decode_T_289; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_291 = _Inst_decode_T_53 ? 7'h44 : _Inst_decode_T_290; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_292 = _Inst_decode_T_51 ? 7'h73 : _Inst_decode_T_291; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_293 = _Inst_decode_T_49 ? 7'h6a : _Inst_decode_T_292; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_294 = _Inst_decode_T_47 ? 7'h71 : _Inst_decode_T_293; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_295 = _Inst_decode_T_45 ? 7'h40 : _Inst_decode_T_294; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_296 = _Inst_decode_T_43 ? 7'h69 : _Inst_decode_T_295; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_297 = _Inst_decode_T_41 ? 7'h68 : _Inst_decode_T_296; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_298 = _Inst_decode_T_39 ? 7'h11 : _Inst_decode_T_297; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_299 = _Inst_decode_T_37 ? 7'h2 : _Inst_decode_T_298; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_300 = _Inst_decode_T_35 ? 7'h8 : _Inst_decode_T_299; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_301 = _Inst_decode_T_33 ? 7'h6 : _Inst_decode_T_300; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_302 = _Inst_decode_T_31 ? 7'h5 : _Inst_decode_T_301; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_303 = _Inst_decode_T_29 ? 7'h4 : _Inst_decode_T_302; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_304 = _Inst_decode_T_27 ? 7'h3 : _Inst_decode_T_303; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_305 = _Inst_decode_T_25 ? 7'h75 : _Inst_decode_T_304; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_306 = _Inst_decode_T_23 ? 7'h71 : _Inst_decode_T_305; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_307 = _Inst_decode_T_21 ? 7'h72 : _Inst_decode_T_306; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_308 = _Inst_decode_T_19 ? 7'he : _Inst_decode_T_307; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_309 = _Inst_decode_T_17 ? 7'h6f : _Inst_decode_T_308; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_310 = _Inst_decode_T_15 ? 7'h6e : _Inst_decode_T_309; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_311 = _Inst_decode_T_13 ? 7'h6d : _Inst_decode_T_310; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_312 = _Inst_decode_T_11 ? 7'h6a : _Inst_decode_T_311; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_313 = _Inst_decode_T_9 ? 7'h47 : _Inst_decode_T_312; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_314 = _Inst_decode_T_7 ? 7'h45 : _Inst_decode_T_313; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_315 = _Inst_decode_T_5 ? 7'h44 : _Inst_decode_T_314; // @[Lookup.scala 34:39]
  wire [6:0] _Inst_decode_T_316 = _Inst_decode_T_3 ? 7'h41 : _Inst_decode_T_315; // @[Lookup.scala 34:39]
  wire [6:0] Inst_decode_2 = _Inst_decode_T_1 ? 7'h40 : _Inst_decode_T_316; // @[Lookup.scala 34:39]
  wire  _Inst_decode_T_321 = _Inst_decode_T_119 ? 1'h0 : _Inst_decode_T_121 | _Inst_decode_T_123; // @[Lookup.scala 34:39]
  wire  _Inst_decode_T_322 = _Inst_decode_T_117 ? 1'h0 : _Inst_decode_T_321; // @[Lookup.scala 34:39]
  wire  _Inst_decode_T_323 = _Inst_decode_T_115 ? 1'h0 : _Inst_decode_T_322; // @[Lookup.scala 34:39]
  wire  _Inst_decode_T_324 = _Inst_decode_T_113 ? 1'h0 : _Inst_decode_T_323; // @[Lookup.scala 34:39]
  wire  _Inst_decode_T_325 = _Inst_decode_T_111 ? 1'h0 : _Inst_decode_T_324; // @[Lookup.scala 34:39]
  wire  _Inst_decode_T_326 = _Inst_decode_T_109 ? 1'h0 : _Inst_decode_T_325; // @[Lookup.scala 34:39]
  wire  _Inst_decode_T_329 = _Inst_decode_T_103 ? 1'h0 : _Inst_decode_T_105 | (_Inst_decode_T_107 | _Inst_decode_T_326); // @[Lookup.scala 34:39]
  wire  _Inst_decode_T_330 = _Inst_decode_T_101 ? 1'h0 : _Inst_decode_T_329; // @[Lookup.scala 34:39]
  wire  _Inst_decode_T_331 = _Inst_decode_T_99 ? 1'h0 : _Inst_decode_T_330; // @[Lookup.scala 34:39]
  wire  _Inst_decode_T_332 = _Inst_decode_T_97 ? 1'h0 : _Inst_decode_T_331; // @[Lookup.scala 34:39]
  wire  _Inst_decode_T_333 = _Inst_decode_T_95 ? 1'h0 : _Inst_decode_T_332; // @[Lookup.scala 34:39]
  wire  _Inst_decode_T_363 = _Inst_decode_T_35 | (_Inst_decode_T_37 | (_Inst_decode_T_39 | (_Inst_decode_T_41 | (
    _Inst_decode_T_43 | (_Inst_decode_T_45 | (_Inst_decode_T_47 | (_Inst_decode_T_49 | (_Inst_decode_T_51 | (
    _Inst_decode_T_53 | (_Inst_decode_T_55 | (_Inst_decode_T_57 | (_Inst_decode_T_59 | (_Inst_decode_T_61 | (
    _Inst_decode_T_63 | (_Inst_decode_T_65 | (_Inst_decode_T_67 | (_Inst_decode_T_69 | (_Inst_decode_T_71 | (
    _Inst_decode_T_73 | (_Inst_decode_T_75 | (_Inst_decode_T_77 | (_Inst_decode_T_79 | (_Inst_decode_T_81 | (
    _Inst_decode_T_83 | (_Inst_decode_T_85 | (_Inst_decode_T_87 | (_Inst_decode_T_89 | (_Inst_decode_T_91 | (
    _Inst_decode_T_93 | _Inst_decode_T_333))))))))))))))))))))))))))))); // @[Lookup.scala 34:39]
  wire  Inst_decode_3 = _Inst_decode_T_1 | (_Inst_decode_T_3 | (_Inst_decode_T_5 | (_Inst_decode_T_7 | (_Inst_decode_T_9
     | (_Inst_decode_T_11 | (_Inst_decode_T_13 | (_Inst_decode_T_15 | (_Inst_decode_T_17 | (_Inst_decode_T_19 | (
    _Inst_decode_T_21 | (_Inst_decode_T_23 | (_Inst_decode_T_25 | (_Inst_decode_T_27 | (_Inst_decode_T_29 | (
    _Inst_decode_T_31 | (_Inst_decode_T_33 | _Inst_decode_T_363)))))))))))))))); // @[Lookup.scala 34:39]
  wire  _srctype1_T = 4'h8 == Inst_decode_0; // @[util.scala 45:32]
  wire  _srctype1_T_2 = 4'h9 == Inst_decode_0; // @[util.scala 45:32]
  wire  _srctype1_T_3 = 4'hb == Inst_decode_0; // @[util.scala 45:32]
  wire  _srctype1_T_4 = 4'h7 == Inst_decode_0; // @[util.scala 45:32]
  wire  _srctype1_T_5 = 4'h3 == Inst_decode_0; // @[util.scala 45:32]
  wire [1:0] _srctype1_T_11 = _srctype1_T_4 ? 2'h2 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _srctype1_T_12 = _srctype1_T_5 ? 2'h2 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] srctype1 = _srctype1_T_11 | _srctype1_T_12; // @[Mux.scala 27:73]
  wire  srctype2 = _srctype1_T | _srctype1_T_4 | _srctype1_T_5; // @[Mux.scala 27:73]
  wire  sign = io_in_bits_Inst[31]; // @[util.scala 11:19]
  wire [51:0] _T_2 = sign ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _T_3 = {_T_2,io_in_bits_Inst[31:20]}; // @[Cat.scala 31:58]
  wire [19:0] _T_7 = {io_in_bits_Inst[19:12],io_in_bits_Inst[20],io_in_bits_Inst[30:21],1'h0}; // @[Cat.scala 31:58]
  wire  sign_1 = _T_7[19]; // @[util.scala 11:19]
  wire [43:0] _T_9 = sign_1 ? 44'hfffffffffff : 44'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _T_10 = {_T_9,io_in_bits_Inst[19:12],io_in_bits_Inst[20],io_in_bits_Inst[30:21],1'h0}; // @[Cat.scala 31:58]
  wire [31:0] _T_13 = {io_in_bits_Inst[31:12],12'h0}; // @[Cat.scala 31:58]
  wire  sign_2 = _T_13[31]; // @[util.scala 11:19]
  wire [31:0] _T_15 = sign_2 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _T_16 = {_T_15,io_in_bits_Inst[31:12],12'h0}; // @[Cat.scala 31:58]
  wire [11:0] _T_19 = {io_in_bits_Inst[31:25],rd}; // @[Cat.scala 31:58]
  wire  sign_3 = _T_19[11]; // @[util.scala 11:19]
  wire [51:0] _T_21 = sign_3 ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _T_22 = {_T_21,io_in_bits_Inst[31:25],rd}; // @[Cat.scala 31:58]
  wire [12:0] _T_27 = {io_in_bits_Inst[31],io_in_bits_Inst[7],io_in_bits_Inst[30:25],io_in_bits_Inst[11:8],1'h0}; // @[Cat.scala 31:58]
  wire  sign_4 = _T_27[12]; // @[util.scala 11:19]
  wire [50:0] _T_29 = sign_4 ? 51'h7ffffffffffff : 51'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _T_30 = {_T_29,io_in_bits_Inst[31],io_in_bits_Inst[7],io_in_bits_Inst[30:25],io_in_bits_Inst[11:8],1'h0}; // @[Cat.scala 31:58]
  wire [63:0] _imm_T_5 = _srctype1_T ? _T_3 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _imm_T_6 = _srctype1_T_4 ? _T_10 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _imm_T_7 = _srctype1_T_5 ? _T_16 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _imm_T_8 = _srctype1_T_2 ? _T_22 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _imm_T_9 = _srctype1_T_3 ? _T_30 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _imm_T_10 = _imm_T_5 | _imm_T_6; // @[Mux.scala 27:73]
  wire [63:0] _imm_T_11 = _imm_T_10 | _imm_T_7; // @[Mux.scala 27:73]
  wire [63:0] _imm_T_12 = _imm_T_11 | _imm_T_8; // @[Mux.scala 27:73]
  assign io_in_ready = io_out_ready; // @[ID.scala 106:15]
  assign io_out_valid = io_in_valid; // @[ID.scala 105:22]
  assign io_out_bits_ctrl_signal_src1Type = {{1'd0}, srctype1}; // @[ID.scala 87:36]
  assign io_out_bits_ctrl_signal_src2Type = {{2'd0}, srctype2}; // @[ID.scala 88:36]
  assign io_out_bits_ctrl_signal_fuType = _Inst_decode_T_1 ? 3'h0 : _Inst_decode_T_253; // @[Lookup.scala 34:39]
  assign io_out_bits_ctrl_signal_inst_valid = Inst_decode_2 == 7'h0 | io_flush | ~io_in_valid ? 1'h0 : 1'h1; // @[ID.scala 89:44]
  assign io_out_bits_ctrl_signal_rfSrc1 = io_in_bits_Inst[19:15]; // @[ID.scala 51:38]
  assign io_out_bits_ctrl_signal_rfSrc2 = io_in_bits_Inst[24:20]; // @[ID.scala 51:63]
  assign io_out_bits_ctrl_signal_rfWen = io_in_valid & Inst_decode_3; // @[ID.scala 84:39]
  assign io_out_bits_ctrl_signal_aluoptype = _Inst_decode_T_1 ? 7'h40 : _Inst_decode_T_316; // @[Lookup.scala 34:39]
  assign io_out_bits_ctrl_signal_rfDest = io_in_bits_Inst[11:7]; // @[ID.scala 51:88]
  assign io_out_bits_ctrl_data_src1 = io_REG1; // @[ID.scala 99:30]
  assign io_out_bits_ctrl_data_src2 = io_REG2; // @[ID.scala 100:30]
  assign io_out_bits_ctrl_data_Imm = _imm_T_12 | _imm_T_9; // @[Mux.scala 27:73]
  assign io_out_bits_ctrl_flow_PC = io_in_bits_PC; // @[ID.scala 92:28]
  assign io_out_bits_ctrl_flow_inst = io_in_bits_Inst; // @[ID.scala 93:30]
endmodule
module Improved_Partial_product(
  input  [2:0]  io_y_3,
  input  [65:0] io_x,
  output [65:0] io_p,
  output [1:0]  io_carry
);
  wire  _io_p_T = io_y_3 == 3'h0; // @[MUL.scala 58:13]
  wire  _io_p_T_1 = io_y_3 == 3'h1; // @[MUL.scala 59:13]
  wire  _io_p_T_2 = io_y_3 == 3'h2; // @[MUL.scala 60:13]
  wire  _io_p_T_3 = io_y_3 == 3'h3; // @[MUL.scala 61:13]
  wire [66:0] _io_p_T_4 = {io_x, 1'h0}; // @[MUL.scala 61:36]
  wire  _io_p_T_5 = io_y_3 == 3'h4; // @[MUL.scala 62:13]
  wire [65:0] _io_p_T_6 = ~io_x; // @[MUL.scala 62:32]
  wire [66:0] _io_p_T_7 = {_io_p_T_6, 1'h0}; // @[MUL.scala 62:39]
  wire  _io_p_T_8 = io_y_3 == 3'h5; // @[MUL.scala 63:13]
  wire  _io_p_T_10 = io_y_3 == 3'h6; // @[MUL.scala 64:13]
  wire [65:0] _io_p_T_14 = _io_p_T_10 ? _io_p_T_6 : 66'h0; // @[Mux.scala 101:16]
  wire [65:0] _io_p_T_15 = _io_p_T_8 ? _io_p_T_6 : _io_p_T_14; // @[Mux.scala 101:16]
  wire [66:0] _io_p_T_16 = _io_p_T_5 ? _io_p_T_7 : {{1'd0}, _io_p_T_15}; // @[Mux.scala 101:16]
  wire [66:0] _io_p_T_17 = _io_p_T_3 ? _io_p_T_4 : _io_p_T_16; // @[Mux.scala 101:16]
  wire [66:0] _io_p_T_18 = _io_p_T_2 ? {{1'd0}, io_x} : _io_p_T_17; // @[Mux.scala 101:16]
  wire [66:0] _io_p_T_19 = _io_p_T_1 ? {{1'd0}, io_x} : _io_p_T_18; // @[Mux.scala 101:16]
  wire [66:0] _io_p_T_20 = _io_p_T ? 67'h0 : _io_p_T_19; // @[Mux.scala 101:16]
  wire [1:0] _io_carry_T_9 = _io_p_T_10 ? 2'h1 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _io_carry_T_10 = _io_p_T_8 ? 2'h1 : _io_carry_T_9; // @[Mux.scala 101:16]
  wire [1:0] _io_carry_T_11 = _io_p_T_5 ? 2'h2 : _io_carry_T_10; // @[Mux.scala 101:16]
  wire [1:0] _io_carry_T_12 = _io_p_T_3 ? 2'h0 : _io_carry_T_11; // @[Mux.scala 101:16]
  wire [1:0] _io_carry_T_13 = _io_p_T_2 ? 2'h0 : _io_carry_T_12; // @[Mux.scala 101:16]
  wire [1:0] _io_carry_T_14 = _io_p_T_1 ? 2'h0 : _io_carry_T_13; // @[Mux.scala 101:16]
  assign io_p = _io_p_T_20[65:0]; // @[MUL.scala 57:8]
  assign io_carry = _io_p_T ? 2'h0 : _io_carry_T_14; // @[Mux.scala 101:16]
endmodule
module Half_Adder(
  input   io_in_0,
  input   io_in_1,
  output  io_out_0,
  output  io_out_1
);
  assign io_out_0 = io_in_0 ^ io_in_1; // @[MUL.scala 119:25]
  assign io_out_1 = io_in_0 & io_in_1; // @[MUL.scala 120:25]
endmodule
module Adder(
  input   io_x1,
  input   io_x2,
  input   io_x3,
  output  io_s,
  output  io_cout
);
  assign io_s = io_x1 ^ io_x2 ^ io_x3; // @[MUL.scala 96:25]
  assign io_cout = io_x1 & io_x2 | io_x1 & io_x3 | io_x2 & io_x3; // @[MUL.scala 97:48]
endmodule
module Booth_Walloc_MUL(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [63:0] io_in_bits_ctrl_data_src1,
  input  [63:0] io_in_bits_ctrl_data_src2,
  output        io_out_valid,
  output [63:0] io_out_bits_result_result_lo
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1545;
  reg [31:0] _RAND_1546;
  reg [31:0] _RAND_1547;
  reg [31:0] _RAND_1548;
  reg [31:0] _RAND_1549;
  reg [31:0] _RAND_1550;
  reg [31:0] _RAND_1551;
  reg [31:0] _RAND_1552;
  reg [31:0] _RAND_1553;
  reg [31:0] _RAND_1554;
  reg [31:0] _RAND_1555;
  reg [31:0] _RAND_1556;
  reg [31:0] _RAND_1557;
  reg [31:0] _RAND_1558;
  reg [31:0] _RAND_1559;
  reg [31:0] _RAND_1560;
  reg [31:0] _RAND_1561;
  reg [31:0] _RAND_1562;
  reg [31:0] _RAND_1563;
  reg [31:0] _RAND_1564;
  reg [31:0] _RAND_1565;
  reg [31:0] _RAND_1566;
  reg [31:0] _RAND_1567;
  reg [31:0] _RAND_1568;
  reg [31:0] _RAND_1569;
  reg [31:0] _RAND_1570;
  reg [31:0] _RAND_1571;
  reg [31:0] _RAND_1572;
  reg [31:0] _RAND_1573;
  reg [31:0] _RAND_1574;
  reg [31:0] _RAND_1575;
  reg [31:0] _RAND_1576;
  reg [31:0] _RAND_1577;
  reg [31:0] _RAND_1578;
  reg [31:0] _RAND_1579;
  reg [31:0] _RAND_1580;
  reg [31:0] _RAND_1581;
  reg [31:0] _RAND_1582;
  reg [31:0] _RAND_1583;
  reg [31:0] _RAND_1584;
  reg [31:0] _RAND_1585;
  reg [31:0] _RAND_1586;
  reg [31:0] _RAND_1587;
  reg [31:0] _RAND_1588;
  reg [31:0] _RAND_1589;
  reg [31:0] _RAND_1590;
  reg [31:0] _RAND_1591;
  reg [31:0] _RAND_1592;
  reg [31:0] _RAND_1593;
  reg [31:0] _RAND_1594;
  reg [31:0] _RAND_1595;
  reg [31:0] _RAND_1596;
  reg [31:0] _RAND_1597;
  reg [31:0] _RAND_1598;
  reg [31:0] _RAND_1599;
  reg [31:0] _RAND_1600;
  reg [31:0] _RAND_1601;
  reg [31:0] _RAND_1602;
  reg [31:0] _RAND_1603;
  reg [31:0] _RAND_1604;
  reg [31:0] _RAND_1605;
  reg [31:0] _RAND_1606;
  reg [31:0] _RAND_1607;
  reg [31:0] _RAND_1608;
  reg [31:0] _RAND_1609;
  reg [31:0] _RAND_1610;
  reg [31:0] _RAND_1611;
  reg [31:0] _RAND_1612;
  reg [31:0] _RAND_1613;
  reg [31:0] _RAND_1614;
  reg [31:0] _RAND_1615;
  reg [31:0] _RAND_1616;
  reg [31:0] _RAND_1617;
  reg [31:0] _RAND_1618;
  reg [31:0] _RAND_1619;
  reg [31:0] _RAND_1620;
  reg [31:0] _RAND_1621;
  reg [31:0] _RAND_1622;
  reg [31:0] _RAND_1623;
  reg [31:0] _RAND_1624;
  reg [31:0] _RAND_1625;
  reg [31:0] _RAND_1626;
  reg [31:0] _RAND_1627;
  reg [31:0] _RAND_1628;
  reg [31:0] _RAND_1629;
  reg [31:0] _RAND_1630;
  reg [31:0] _RAND_1631;
  reg [31:0] _RAND_1632;
  reg [31:0] _RAND_1633;
  reg [31:0] _RAND_1634;
  reg [31:0] _RAND_1635;
  reg [31:0] _RAND_1636;
  reg [31:0] _RAND_1637;
  reg [31:0] _RAND_1638;
  reg [31:0] _RAND_1639;
  reg [31:0] _RAND_1640;
  reg [31:0] _RAND_1641;
  reg [31:0] _RAND_1642;
  reg [31:0] _RAND_1643;
  reg [31:0] _RAND_1644;
  reg [31:0] _RAND_1645;
  reg [31:0] _RAND_1646;
  reg [31:0] _RAND_1647;
  reg [31:0] _RAND_1648;
  reg [31:0] _RAND_1649;
  reg [31:0] _RAND_1650;
  reg [31:0] _RAND_1651;
  reg [31:0] _RAND_1652;
  reg [31:0] _RAND_1653;
  reg [31:0] _RAND_1654;
  reg [31:0] _RAND_1655;
  reg [31:0] _RAND_1656;
  reg [31:0] _RAND_1657;
  reg [31:0] _RAND_1658;
  reg [31:0] _RAND_1659;
  reg [31:0] _RAND_1660;
  reg [31:0] _RAND_1661;
  reg [31:0] _RAND_1662;
  reg [31:0] _RAND_1663;
  reg [31:0] _RAND_1664;
  reg [31:0] _RAND_1665;
  reg [31:0] _RAND_1666;
  reg [31:0] _RAND_1667;
  reg [31:0] _RAND_1668;
  reg [31:0] _RAND_1669;
  reg [31:0] _RAND_1670;
  reg [31:0] _RAND_1671;
  reg [31:0] _RAND_1672;
  reg [31:0] _RAND_1673;
  reg [31:0] _RAND_1674;
  reg [31:0] _RAND_1675;
  reg [31:0] _RAND_1676;
  reg [31:0] _RAND_1677;
  reg [31:0] _RAND_1678;
  reg [31:0] _RAND_1679;
  reg [31:0] _RAND_1680;
  reg [31:0] _RAND_1681;
  reg [31:0] _RAND_1682;
  reg [31:0] _RAND_1683;
  reg [31:0] _RAND_1684;
  reg [31:0] _RAND_1685;
  reg [31:0] _RAND_1686;
  reg [31:0] _RAND_1687;
  reg [31:0] _RAND_1688;
  reg [31:0] _RAND_1689;
  reg [31:0] _RAND_1690;
  reg [31:0] _RAND_1691;
  reg [31:0] _RAND_1692;
  reg [31:0] _RAND_1693;
  reg [31:0] _RAND_1694;
  reg [31:0] _RAND_1695;
  reg [31:0] _RAND_1696;
  reg [31:0] _RAND_1697;
  reg [31:0] _RAND_1698;
  reg [31:0] _RAND_1699;
  reg [31:0] _RAND_1700;
  reg [31:0] _RAND_1701;
  reg [31:0] _RAND_1702;
  reg [31:0] _RAND_1703;
  reg [31:0] _RAND_1704;
  reg [31:0] _RAND_1705;
  reg [31:0] _RAND_1706;
  reg [31:0] _RAND_1707;
  reg [31:0] _RAND_1708;
  reg [31:0] _RAND_1709;
  reg [31:0] _RAND_1710;
  reg [31:0] _RAND_1711;
  reg [31:0] _RAND_1712;
  reg [31:0] _RAND_1713;
  reg [31:0] _RAND_1714;
  reg [31:0] _RAND_1715;
  reg [31:0] _RAND_1716;
  reg [31:0] _RAND_1717;
  reg [31:0] _RAND_1718;
  reg [31:0] _RAND_1719;
  reg [31:0] _RAND_1720;
  reg [31:0] _RAND_1721;
  reg [31:0] _RAND_1722;
  reg [31:0] _RAND_1723;
  reg [31:0] _RAND_1724;
  reg [31:0] _RAND_1725;
  reg [31:0] _RAND_1726;
  reg [31:0] _RAND_1727;
  reg [31:0] _RAND_1728;
  reg [31:0] _RAND_1729;
  reg [31:0] _RAND_1730;
  reg [31:0] _RAND_1731;
  reg [31:0] _RAND_1732;
  reg [31:0] _RAND_1733;
  reg [31:0] _RAND_1734;
  reg [31:0] _RAND_1735;
  reg [31:0] _RAND_1736;
  reg [31:0] _RAND_1737;
  reg [31:0] _RAND_1738;
  reg [31:0] _RAND_1739;
  reg [31:0] _RAND_1740;
  reg [31:0] _RAND_1741;
  reg [31:0] _RAND_1742;
  reg [31:0] _RAND_1743;
  reg [31:0] _RAND_1744;
  reg [31:0] _RAND_1745;
  reg [31:0] _RAND_1746;
  reg [31:0] _RAND_1747;
  reg [31:0] _RAND_1748;
  reg [31:0] _RAND_1749;
  reg [31:0] _RAND_1750;
  reg [31:0] _RAND_1751;
  reg [31:0] _RAND_1752;
  reg [31:0] _RAND_1753;
  reg [31:0] _RAND_1754;
  reg [31:0] _RAND_1755;
  reg [31:0] _RAND_1756;
  reg [31:0] _RAND_1757;
  reg [31:0] _RAND_1758;
  reg [31:0] _RAND_1759;
  reg [31:0] _RAND_1760;
  reg [31:0] _RAND_1761;
  reg [31:0] _RAND_1762;
  reg [31:0] _RAND_1763;
  reg [31:0] _RAND_1764;
  reg [31:0] _RAND_1765;
  reg [31:0] _RAND_1766;
  reg [31:0] _RAND_1767;
  reg [31:0] _RAND_1768;
  reg [31:0] _RAND_1769;
  reg [31:0] _RAND_1770;
  reg [31:0] _RAND_1771;
  reg [31:0] _RAND_1772;
  reg [31:0] _RAND_1773;
  reg [31:0] _RAND_1774;
  reg [31:0] _RAND_1775;
  reg [31:0] _RAND_1776;
  reg [31:0] _RAND_1777;
  reg [31:0] _RAND_1778;
  reg [31:0] _RAND_1779;
  reg [31:0] _RAND_1780;
  reg [31:0] _RAND_1781;
  reg [31:0] _RAND_1782;
  reg [31:0] _RAND_1783;
  reg [31:0] _RAND_1784;
  reg [31:0] _RAND_1785;
  reg [31:0] _RAND_1786;
  reg [31:0] _RAND_1787;
  reg [31:0] _RAND_1788;
  reg [31:0] _RAND_1789;
  reg [31:0] _RAND_1790;
  reg [31:0] _RAND_1791;
  reg [31:0] _RAND_1792;
  reg [31:0] _RAND_1793;
  reg [31:0] _RAND_1794;
  reg [31:0] _RAND_1795;
  reg [31:0] _RAND_1796;
  reg [31:0] _RAND_1797;
  reg [31:0] _RAND_1798;
  reg [31:0] _RAND_1799;
  reg [31:0] _RAND_1800;
  reg [31:0] _RAND_1801;
  reg [31:0] _RAND_1802;
  reg [31:0] _RAND_1803;
  reg [31:0] _RAND_1804;
  reg [31:0] _RAND_1805;
  reg [31:0] _RAND_1806;
  reg [31:0] _RAND_1807;
  reg [31:0] _RAND_1808;
  reg [31:0] _RAND_1809;
  reg [31:0] _RAND_1810;
  reg [31:0] _RAND_1811;
  reg [31:0] _RAND_1812;
  reg [31:0] _RAND_1813;
  reg [31:0] _RAND_1814;
  reg [31:0] _RAND_1815;
  reg [31:0] _RAND_1816;
  reg [31:0] _RAND_1817;
  reg [31:0] _RAND_1818;
  reg [31:0] _RAND_1819;
  reg [31:0] _RAND_1820;
  reg [31:0] _RAND_1821;
  reg [31:0] _RAND_1822;
  reg [31:0] _RAND_1823;
  reg [31:0] _RAND_1824;
  reg [31:0] _RAND_1825;
  reg [31:0] _RAND_1826;
  reg [31:0] _RAND_1827;
  reg [31:0] _RAND_1828;
  reg [31:0] _RAND_1829;
  reg [31:0] _RAND_1830;
  reg [31:0] _RAND_1831;
  reg [31:0] _RAND_1832;
  reg [31:0] _RAND_1833;
  reg [31:0] _RAND_1834;
  reg [31:0] _RAND_1835;
  reg [31:0] _RAND_1836;
  reg [31:0] _RAND_1837;
  reg [31:0] _RAND_1838;
  reg [31:0] _RAND_1839;
  reg [31:0] _RAND_1840;
  reg [31:0] _RAND_1841;
  reg [31:0] _RAND_1842;
  reg [31:0] _RAND_1843;
  reg [31:0] _RAND_1844;
  reg [31:0] _RAND_1845;
  reg [31:0] _RAND_1846;
  reg [31:0] _RAND_1847;
  reg [31:0] _RAND_1848;
  reg [31:0] _RAND_1849;
  reg [31:0] _RAND_1850;
  reg [31:0] _RAND_1851;
  reg [31:0] _RAND_1852;
  reg [31:0] _RAND_1853;
  reg [31:0] _RAND_1854;
  reg [31:0] _RAND_1855;
  reg [31:0] _RAND_1856;
  reg [31:0] _RAND_1857;
  reg [31:0] _RAND_1858;
  reg [31:0] _RAND_1859;
  reg [31:0] _RAND_1860;
  reg [31:0] _RAND_1861;
  reg [31:0] _RAND_1862;
  reg [31:0] _RAND_1863;
  reg [31:0] _RAND_1864;
  reg [31:0] _RAND_1865;
  reg [31:0] _RAND_1866;
  reg [31:0] _RAND_1867;
  reg [31:0] _RAND_1868;
  reg [31:0] _RAND_1869;
  reg [31:0] _RAND_1870;
  reg [31:0] _RAND_1871;
  reg [31:0] _RAND_1872;
  reg [31:0] _RAND_1873;
  reg [31:0] _RAND_1874;
  reg [31:0] _RAND_1875;
  reg [31:0] _RAND_1876;
  reg [31:0] _RAND_1877;
  reg [31:0] _RAND_1878;
  reg [31:0] _RAND_1879;
  reg [31:0] _RAND_1880;
  reg [31:0] _RAND_1881;
  reg [31:0] _RAND_1882;
  reg [31:0] _RAND_1883;
  reg [31:0] _RAND_1884;
  reg [31:0] _RAND_1885;
  reg [31:0] _RAND_1886;
  reg [31:0] _RAND_1887;
  reg [31:0] _RAND_1888;
  reg [31:0] _RAND_1889;
  reg [31:0] _RAND_1890;
  reg [31:0] _RAND_1891;
  reg [31:0] _RAND_1892;
  reg [31:0] _RAND_1893;
  reg [31:0] _RAND_1894;
  reg [31:0] _RAND_1895;
  reg [31:0] _RAND_1896;
  reg [31:0] _RAND_1897;
  reg [31:0] _RAND_1898;
  reg [31:0] _RAND_1899;
  reg [31:0] _RAND_1900;
  reg [31:0] _RAND_1901;
  reg [31:0] _RAND_1902;
  reg [31:0] _RAND_1903;
  reg [31:0] _RAND_1904;
  reg [31:0] _RAND_1905;
  reg [31:0] _RAND_1906;
  reg [31:0] _RAND_1907;
  reg [31:0] _RAND_1908;
  reg [31:0] _RAND_1909;
  reg [31:0] _RAND_1910;
  reg [31:0] _RAND_1911;
  reg [31:0] _RAND_1912;
  reg [31:0] _RAND_1913;
  reg [31:0] _RAND_1914;
  reg [31:0] _RAND_1915;
  reg [31:0] _RAND_1916;
  reg [31:0] _RAND_1917;
  reg [31:0] _RAND_1918;
  reg [31:0] _RAND_1919;
  reg [31:0] _RAND_1920;
  reg [31:0] _RAND_1921;
  reg [31:0] _RAND_1922;
  reg [31:0] _RAND_1923;
  reg [31:0] _RAND_1924;
  reg [31:0] _RAND_1925;
  reg [31:0] _RAND_1926;
  reg [31:0] _RAND_1927;
  reg [31:0] _RAND_1928;
  reg [31:0] _RAND_1929;
  reg [31:0] _RAND_1930;
  reg [31:0] _RAND_1931;
  reg [31:0] _RAND_1932;
  reg [31:0] _RAND_1933;
  reg [31:0] _RAND_1934;
  reg [31:0] _RAND_1935;
  reg [31:0] _RAND_1936;
  reg [31:0] _RAND_1937;
  reg [31:0] _RAND_1938;
  reg [31:0] _RAND_1939;
  reg [31:0] _RAND_1940;
  reg [31:0] _RAND_1941;
  reg [31:0] _RAND_1942;
  reg [31:0] _RAND_1943;
  reg [31:0] _RAND_1944;
  reg [31:0] _RAND_1945;
  reg [31:0] _RAND_1946;
  reg [31:0] _RAND_1947;
  reg [31:0] _RAND_1948;
  reg [31:0] _RAND_1949;
  reg [31:0] _RAND_1950;
  reg [31:0] _RAND_1951;
  reg [31:0] _RAND_1952;
  reg [31:0] _RAND_1953;
  reg [31:0] _RAND_1954;
  reg [31:0] _RAND_1955;
  reg [31:0] _RAND_1956;
  reg [31:0] _RAND_1957;
  reg [31:0] _RAND_1958;
  reg [31:0] _RAND_1959;
  reg [31:0] _RAND_1960;
  reg [31:0] _RAND_1961;
  reg [31:0] _RAND_1962;
  reg [31:0] _RAND_1963;
  reg [31:0] _RAND_1964;
  reg [31:0] _RAND_1965;
  reg [31:0] _RAND_1966;
  reg [31:0] _RAND_1967;
  reg [31:0] _RAND_1968;
  reg [31:0] _RAND_1969;
  reg [31:0] _RAND_1970;
  reg [31:0] _RAND_1971;
  reg [31:0] _RAND_1972;
  reg [31:0] _RAND_1973;
  reg [31:0] _RAND_1974;
  reg [31:0] _RAND_1975;
  reg [31:0] _RAND_1976;
  reg [31:0] _RAND_1977;
  reg [31:0] _RAND_1978;
  reg [31:0] _RAND_1979;
  reg [31:0] _RAND_1980;
  reg [31:0] _RAND_1981;
  reg [31:0] _RAND_1982;
  reg [31:0] _RAND_1983;
  reg [31:0] _RAND_1984;
  reg [31:0] _RAND_1985;
  reg [31:0] _RAND_1986;
  reg [31:0] _RAND_1987;
  reg [31:0] _RAND_1988;
  reg [31:0] _RAND_1989;
  reg [31:0] _RAND_1990;
  reg [31:0] _RAND_1991;
  reg [31:0] _RAND_1992;
  reg [31:0] _RAND_1993;
  reg [31:0] _RAND_1994;
  reg [31:0] _RAND_1995;
  reg [31:0] _RAND_1996;
  reg [31:0] _RAND_1997;
  reg [31:0] _RAND_1998;
  reg [31:0] _RAND_1999;
  reg [31:0] _RAND_2000;
  reg [31:0] _RAND_2001;
  reg [31:0] _RAND_2002;
  reg [31:0] _RAND_2003;
  reg [31:0] _RAND_2004;
  reg [31:0] _RAND_2005;
  reg [31:0] _RAND_2006;
  reg [31:0] _RAND_2007;
  reg [31:0] _RAND_2008;
  reg [31:0] _RAND_2009;
  reg [31:0] _RAND_2010;
  reg [31:0] _RAND_2011;
  reg [31:0] _RAND_2012;
  reg [31:0] _RAND_2013;
  reg [31:0] _RAND_2014;
  reg [31:0] _RAND_2015;
  reg [31:0] _RAND_2016;
  reg [31:0] _RAND_2017;
  reg [31:0] _RAND_2018;
  reg [31:0] _RAND_2019;
  reg [31:0] _RAND_2020;
  reg [31:0] _RAND_2021;
  reg [31:0] _RAND_2022;
  reg [31:0] _RAND_2023;
  reg [31:0] _RAND_2024;
  reg [31:0] _RAND_2025;
  reg [31:0] _RAND_2026;
  reg [31:0] _RAND_2027;
  reg [31:0] _RAND_2028;
  reg [31:0] _RAND_2029;
  reg [31:0] _RAND_2030;
  reg [31:0] _RAND_2031;
  reg [31:0] _RAND_2032;
  reg [31:0] _RAND_2033;
  reg [31:0] _RAND_2034;
  reg [31:0] _RAND_2035;
  reg [31:0] _RAND_2036;
  reg [31:0] _RAND_2037;
  reg [31:0] _RAND_2038;
  reg [31:0] _RAND_2039;
  reg [31:0] _RAND_2040;
  reg [31:0] _RAND_2041;
  reg [31:0] _RAND_2042;
  reg [31:0] _RAND_2043;
  reg [31:0] _RAND_2044;
  reg [31:0] _RAND_2045;
  reg [31:0] _RAND_2046;
  reg [31:0] _RAND_2047;
  reg [31:0] _RAND_2048;
  reg [31:0] _RAND_2049;
  reg [31:0] _RAND_2050;
  reg [31:0] _RAND_2051;
  reg [31:0] _RAND_2052;
  reg [31:0] _RAND_2053;
  reg [31:0] _RAND_2054;
  reg [31:0] _RAND_2055;
  reg [31:0] _RAND_2056;
  reg [31:0] _RAND_2057;
  reg [31:0] _RAND_2058;
  reg [31:0] _RAND_2059;
  reg [31:0] _RAND_2060;
  reg [31:0] _RAND_2061;
  reg [31:0] _RAND_2062;
  reg [31:0] _RAND_2063;
  reg [31:0] _RAND_2064;
  reg [31:0] _RAND_2065;
  reg [31:0] _RAND_2066;
  reg [31:0] _RAND_2067;
  reg [31:0] _RAND_2068;
  reg [31:0] _RAND_2069;
  reg [31:0] _RAND_2070;
  reg [31:0] _RAND_2071;
  reg [31:0] _RAND_2072;
  reg [31:0] _RAND_2073;
  reg [31:0] _RAND_2074;
  reg [31:0] _RAND_2075;
  reg [31:0] _RAND_2076;
  reg [31:0] _RAND_2077;
  reg [31:0] _RAND_2078;
  reg [31:0] _RAND_2079;
  reg [31:0] _RAND_2080;
  reg [31:0] _RAND_2081;
  reg [31:0] _RAND_2082;
  reg [31:0] _RAND_2083;
  reg [31:0] _RAND_2084;
  reg [31:0] _RAND_2085;
  reg [31:0] _RAND_2086;
  reg [31:0] _RAND_2087;
  reg [31:0] _RAND_2088;
  reg [31:0] _RAND_2089;
  reg [31:0] _RAND_2090;
  reg [31:0] _RAND_2091;
  reg [31:0] _RAND_2092;
  reg [31:0] _RAND_2093;
  reg [31:0] _RAND_2094;
  reg [31:0] _RAND_2095;
  reg [31:0] _RAND_2096;
  reg [31:0] _RAND_2097;
  reg [31:0] _RAND_2098;
  reg [31:0] _RAND_2099;
  reg [31:0] _RAND_2100;
  reg [31:0] _RAND_2101;
  reg [31:0] _RAND_2102;
  reg [31:0] _RAND_2103;
  reg [31:0] _RAND_2104;
  reg [31:0] _RAND_2105;
  reg [31:0] _RAND_2106;
  reg [31:0] _RAND_2107;
  reg [31:0] _RAND_2108;
  reg [31:0] _RAND_2109;
  reg [31:0] _RAND_2110;
  reg [31:0] _RAND_2111;
  reg [31:0] _RAND_2112;
  reg [31:0] _RAND_2113;
  reg [31:0] _RAND_2114;
  reg [31:0] _RAND_2115;
  reg [31:0] _RAND_2116;
  reg [31:0] _RAND_2117;
  reg [31:0] _RAND_2118;
  reg [31:0] _RAND_2119;
  reg [31:0] _RAND_2120;
  reg [31:0] _RAND_2121;
  reg [31:0] _RAND_2122;
  reg [31:0] _RAND_2123;
  reg [31:0] _RAND_2124;
  reg [31:0] _RAND_2125;
  reg [31:0] _RAND_2126;
  reg [31:0] _RAND_2127;
  reg [31:0] _RAND_2128;
  reg [31:0] _RAND_2129;
  reg [31:0] _RAND_2130;
  reg [31:0] _RAND_2131;
  reg [31:0] _RAND_2132;
  reg [31:0] _RAND_2133;
  reg [31:0] _RAND_2134;
  reg [31:0] _RAND_2135;
  reg [31:0] _RAND_2136;
  reg [31:0] _RAND_2137;
  reg [31:0] _RAND_2138;
  reg [31:0] _RAND_2139;
  reg [31:0] _RAND_2140;
  reg [31:0] _RAND_2141;
  reg [31:0] _RAND_2142;
  reg [31:0] _RAND_2143;
  reg [31:0] _RAND_2144;
  reg [31:0] _RAND_2145;
  reg [31:0] _RAND_2146;
  reg [31:0] _RAND_2147;
  reg [31:0] _RAND_2148;
  reg [31:0] _RAND_2149;
  reg [31:0] _RAND_2150;
  reg [31:0] _RAND_2151;
  reg [31:0] _RAND_2152;
  reg [31:0] _RAND_2153;
  reg [31:0] _RAND_2154;
  reg [31:0] _RAND_2155;
  reg [31:0] _RAND_2156;
  reg [31:0] _RAND_2157;
  reg [31:0] _RAND_2158;
  reg [31:0] _RAND_2159;
  reg [31:0] _RAND_2160;
  reg [31:0] _RAND_2161;
  reg [31:0] _RAND_2162;
  reg [31:0] _RAND_2163;
  reg [31:0] _RAND_2164;
  reg [31:0] _RAND_2165;
  reg [31:0] _RAND_2166;
  reg [31:0] _RAND_2167;
  reg [31:0] _RAND_2168;
  reg [31:0] _RAND_2169;
  reg [31:0] _RAND_2170;
  reg [31:0] _RAND_2171;
  reg [31:0] _RAND_2172;
  reg [31:0] _RAND_2173;
  reg [31:0] _RAND_2174;
  reg [31:0] _RAND_2175;
  reg [31:0] _RAND_2176;
  reg [31:0] _RAND_2177;
  reg [31:0] _RAND_2178;
  reg [31:0] _RAND_2179;
  reg [31:0] _RAND_2180;
  reg [31:0] _RAND_2181;
  reg [31:0] _RAND_2182;
  reg [31:0] _RAND_2183;
  reg [31:0] _RAND_2184;
  reg [31:0] _RAND_2185;
  reg [31:0] _RAND_2186;
  reg [31:0] _RAND_2187;
  reg [31:0] _RAND_2188;
  reg [31:0] _RAND_2189;
  reg [31:0] _RAND_2190;
  reg [31:0] _RAND_2191;
  reg [31:0] _RAND_2192;
  reg [31:0] _RAND_2193;
  reg [31:0] _RAND_2194;
  reg [31:0] _RAND_2195;
  reg [31:0] _RAND_2196;
  reg [31:0] _RAND_2197;
  reg [31:0] _RAND_2198;
  reg [31:0] _RAND_2199;
  reg [31:0] _RAND_2200;
  reg [31:0] _RAND_2201;
  reg [31:0] _RAND_2202;
  reg [31:0] _RAND_2203;
  reg [31:0] _RAND_2204;
  reg [31:0] _RAND_2205;
  reg [31:0] _RAND_2206;
  reg [31:0] _RAND_2207;
  reg [31:0] _RAND_2208;
  reg [31:0] _RAND_2209;
  reg [31:0] _RAND_2210;
  reg [31:0] _RAND_2211;
  reg [31:0] _RAND_2212;
  reg [31:0] _RAND_2213;
  reg [31:0] _RAND_2214;
  reg [31:0] _RAND_2215;
  reg [31:0] _RAND_2216;
  reg [31:0] _RAND_2217;
  reg [31:0] _RAND_2218;
  reg [31:0] _RAND_2219;
  reg [31:0] _RAND_2220;
  reg [31:0] _RAND_2221;
  reg [31:0] _RAND_2222;
  reg [31:0] _RAND_2223;
  reg [31:0] _RAND_2224;
  reg [31:0] _RAND_2225;
  reg [31:0] _RAND_2226;
  reg [31:0] _RAND_2227;
  reg [31:0] _RAND_2228;
  reg [31:0] _RAND_2229;
  reg [31:0] _RAND_2230;
  reg [31:0] _RAND_2231;
  reg [31:0] _RAND_2232;
  reg [31:0] _RAND_2233;
  reg [31:0] _RAND_2234;
  reg [31:0] _RAND_2235;
  reg [31:0] _RAND_2236;
  reg [31:0] _RAND_2237;
  reg [31:0] _RAND_2238;
  reg [31:0] _RAND_2239;
  reg [31:0] _RAND_2240;
  reg [31:0] _RAND_2241;
  reg [31:0] _RAND_2242;
  reg [31:0] _RAND_2243;
  reg [31:0] _RAND_2244;
  reg [31:0] _RAND_2245;
  reg [31:0] _RAND_2246;
  reg [31:0] _RAND_2247;
  reg [31:0] _RAND_2248;
  reg [31:0] _RAND_2249;
  reg [31:0] _RAND_2250;
  reg [31:0] _RAND_2251;
  reg [31:0] _RAND_2252;
  reg [31:0] _RAND_2253;
  reg [31:0] _RAND_2254;
  reg [31:0] _RAND_2255;
  reg [31:0] _RAND_2256;
  reg [31:0] _RAND_2257;
  reg [31:0] _RAND_2258;
  reg [31:0] _RAND_2259;
  reg [31:0] _RAND_2260;
  reg [31:0] _RAND_2261;
  reg [31:0] _RAND_2262;
  reg [31:0] _RAND_2263;
  reg [31:0] _RAND_2264;
  reg [31:0] _RAND_2265;
  reg [31:0] _RAND_2266;
  reg [31:0] _RAND_2267;
  reg [31:0] _RAND_2268;
  reg [31:0] _RAND_2269;
  reg [31:0] _RAND_2270;
  reg [31:0] _RAND_2271;
  reg [31:0] _RAND_2272;
  reg [31:0] _RAND_2273;
  reg [31:0] _RAND_2274;
  reg [31:0] _RAND_2275;
  reg [31:0] _RAND_2276;
  reg [31:0] _RAND_2277;
  reg [31:0] _RAND_2278;
  reg [31:0] _RAND_2279;
  reg [31:0] _RAND_2280;
  reg [31:0] _RAND_2281;
  reg [31:0] _RAND_2282;
  reg [31:0] _RAND_2283;
  reg [31:0] _RAND_2284;
  reg [31:0] _RAND_2285;
  reg [31:0] _RAND_2286;
  reg [31:0] _RAND_2287;
  reg [31:0] _RAND_2288;
  reg [31:0] _RAND_2289;
  reg [31:0] _RAND_2290;
  reg [31:0] _RAND_2291;
  reg [31:0] _RAND_2292;
  reg [31:0] _RAND_2293;
  reg [31:0] _RAND_2294;
  reg [31:0] _RAND_2295;
  reg [31:0] _RAND_2296;
  reg [31:0] _RAND_2297;
  reg [31:0] _RAND_2298;
  reg [31:0] _RAND_2299;
  reg [31:0] _RAND_2300;
  reg [31:0] _RAND_2301;
  reg [31:0] _RAND_2302;
  reg [31:0] _RAND_2303;
  reg [31:0] _RAND_2304;
  reg [31:0] _RAND_2305;
  reg [31:0] _RAND_2306;
  reg [31:0] _RAND_2307;
  reg [31:0] _RAND_2308;
  reg [31:0] _RAND_2309;
  reg [31:0] _RAND_2310;
  reg [31:0] _RAND_2311;
  reg [31:0] _RAND_2312;
  reg [31:0] _RAND_2313;
  reg [31:0] _RAND_2314;
  reg [31:0] _RAND_2315;
  reg [31:0] _RAND_2316;
  reg [31:0] _RAND_2317;
  reg [31:0] _RAND_2318;
  reg [31:0] _RAND_2319;
  reg [31:0] _RAND_2320;
  reg [31:0] _RAND_2321;
  reg [31:0] _RAND_2322;
  reg [31:0] _RAND_2323;
  reg [31:0] _RAND_2324;
  reg [31:0] _RAND_2325;
  reg [31:0] _RAND_2326;
  reg [31:0] _RAND_2327;
  reg [31:0] _RAND_2328;
  reg [31:0] _RAND_2329;
  reg [31:0] _RAND_2330;
  reg [31:0] _RAND_2331;
  reg [31:0] _RAND_2332;
  reg [31:0] _RAND_2333;
  reg [31:0] _RAND_2334;
  reg [31:0] _RAND_2335;
  reg [31:0] _RAND_2336;
  reg [31:0] _RAND_2337;
  reg [31:0] _RAND_2338;
  reg [31:0] _RAND_2339;
  reg [31:0] _RAND_2340;
  reg [31:0] _RAND_2341;
  reg [31:0] _RAND_2342;
  reg [31:0] _RAND_2343;
  reg [31:0] _RAND_2344;
  reg [31:0] _RAND_2345;
  reg [31:0] _RAND_2346;
  reg [31:0] _RAND_2347;
  reg [31:0] _RAND_2348;
  reg [31:0] _RAND_2349;
  reg [31:0] _RAND_2350;
  reg [31:0] _RAND_2351;
  reg [31:0] _RAND_2352;
  reg [31:0] _RAND_2353;
  reg [31:0] _RAND_2354;
  reg [31:0] _RAND_2355;
  reg [31:0] _RAND_2356;
  reg [31:0] _RAND_2357;
  reg [31:0] _RAND_2358;
  reg [31:0] _RAND_2359;
  reg [31:0] _RAND_2360;
  reg [31:0] _RAND_2361;
  reg [31:0] _RAND_2362;
  reg [31:0] _RAND_2363;
  reg [31:0] _RAND_2364;
  reg [31:0] _RAND_2365;
  reg [31:0] _RAND_2366;
  reg [31:0] _RAND_2367;
  reg [31:0] _RAND_2368;
  reg [31:0] _RAND_2369;
  reg [31:0] _RAND_2370;
  reg [31:0] _RAND_2371;
  reg [31:0] _RAND_2372;
  reg [31:0] _RAND_2373;
  reg [31:0] _RAND_2374;
  reg [31:0] _RAND_2375;
  reg [31:0] _RAND_2376;
  reg [31:0] _RAND_2377;
  reg [31:0] _RAND_2378;
  reg [31:0] _RAND_2379;
  reg [31:0] _RAND_2380;
  reg [31:0] _RAND_2381;
  reg [31:0] _RAND_2382;
  reg [31:0] _RAND_2383;
  reg [31:0] _RAND_2384;
  reg [31:0] _RAND_2385;
  reg [31:0] _RAND_2386;
  reg [31:0] _RAND_2387;
  reg [31:0] _RAND_2388;
  reg [31:0] _RAND_2389;
  reg [31:0] _RAND_2390;
  reg [31:0] _RAND_2391;
  reg [31:0] _RAND_2392;
  reg [31:0] _RAND_2393;
  reg [31:0] _RAND_2394;
  reg [31:0] _RAND_2395;
  reg [31:0] _RAND_2396;
  reg [31:0] _RAND_2397;
  reg [31:0] _RAND_2398;
  reg [31:0] _RAND_2399;
  reg [31:0] _RAND_2400;
  reg [31:0] _RAND_2401;
  reg [31:0] _RAND_2402;
  reg [31:0] _RAND_2403;
  reg [31:0] _RAND_2404;
  reg [31:0] _RAND_2405;
  reg [31:0] _RAND_2406;
  reg [31:0] _RAND_2407;
  reg [31:0] _RAND_2408;
  reg [31:0] _RAND_2409;
  reg [31:0] _RAND_2410;
  reg [31:0] _RAND_2411;
  reg [31:0] _RAND_2412;
  reg [31:0] _RAND_2413;
  reg [31:0] _RAND_2414;
  reg [31:0] _RAND_2415;
  reg [31:0] _RAND_2416;
  reg [31:0] _RAND_2417;
  reg [31:0] _RAND_2418;
  reg [31:0] _RAND_2419;
  reg [31:0] _RAND_2420;
  reg [31:0] _RAND_2421;
  reg [31:0] _RAND_2422;
  reg [31:0] _RAND_2423;
  reg [31:0] _RAND_2424;
  reg [31:0] _RAND_2425;
  reg [31:0] _RAND_2426;
  reg [31:0] _RAND_2427;
  reg [31:0] _RAND_2428;
  reg [31:0] _RAND_2429;
  reg [31:0] _RAND_2430;
  reg [31:0] _RAND_2431;
  reg [31:0] _RAND_2432;
  reg [31:0] _RAND_2433;
  reg [31:0] _RAND_2434;
  reg [31:0] _RAND_2435;
  reg [31:0] _RAND_2436;
  reg [31:0] _RAND_2437;
  reg [31:0] _RAND_2438;
  reg [31:0] _RAND_2439;
  reg [31:0] _RAND_2440;
  reg [31:0] _RAND_2441;
  reg [31:0] _RAND_2442;
  reg [31:0] _RAND_2443;
  reg [31:0] _RAND_2444;
  reg [31:0] _RAND_2445;
  reg [31:0] _RAND_2446;
  reg [31:0] _RAND_2447;
  reg [31:0] _RAND_2448;
  reg [31:0] _RAND_2449;
  reg [31:0] _RAND_2450;
  reg [31:0] _RAND_2451;
  reg [31:0] _RAND_2452;
  reg [31:0] _RAND_2453;
  reg [31:0] _RAND_2454;
  reg [31:0] _RAND_2455;
  reg [31:0] _RAND_2456;
  reg [31:0] _RAND_2457;
  reg [31:0] _RAND_2458;
  reg [31:0] _RAND_2459;
  reg [31:0] _RAND_2460;
  reg [31:0] _RAND_2461;
  reg [31:0] _RAND_2462;
  reg [31:0] _RAND_2463;
  reg [31:0] _RAND_2464;
  reg [31:0] _RAND_2465;
  reg [31:0] _RAND_2466;
  reg [31:0] _RAND_2467;
  reg [31:0] _RAND_2468;
  reg [31:0] _RAND_2469;
  reg [31:0] _RAND_2470;
  reg [31:0] _RAND_2471;
  reg [31:0] _RAND_2472;
  reg [31:0] _RAND_2473;
  reg [31:0] _RAND_2474;
  reg [31:0] _RAND_2475;
  reg [31:0] _RAND_2476;
  reg [31:0] _RAND_2477;
  reg [31:0] _RAND_2478;
  reg [31:0] _RAND_2479;
  reg [31:0] _RAND_2480;
  reg [31:0] _RAND_2481;
  reg [31:0] _RAND_2482;
  reg [31:0] _RAND_2483;
  reg [31:0] _RAND_2484;
  reg [31:0] _RAND_2485;
  reg [31:0] _RAND_2486;
  reg [31:0] _RAND_2487;
  reg [31:0] _RAND_2488;
  reg [31:0] _RAND_2489;
  reg [31:0] _RAND_2490;
  reg [31:0] _RAND_2491;
  reg [31:0] _RAND_2492;
  reg [31:0] _RAND_2493;
  reg [31:0] _RAND_2494;
  reg [31:0] _RAND_2495;
  reg [31:0] _RAND_2496;
  reg [31:0] _RAND_2497;
  reg [31:0] _RAND_2498;
  reg [31:0] _RAND_2499;
  reg [31:0] _RAND_2500;
  reg [31:0] _RAND_2501;
  reg [31:0] _RAND_2502;
  reg [31:0] _RAND_2503;
  reg [31:0] _RAND_2504;
  reg [31:0] _RAND_2505;
  reg [31:0] _RAND_2506;
  reg [31:0] _RAND_2507;
  reg [31:0] _RAND_2508;
  reg [31:0] _RAND_2509;
  reg [31:0] _RAND_2510;
  reg [31:0] _RAND_2511;
  reg [31:0] _RAND_2512;
  reg [31:0] _RAND_2513;
  reg [31:0] _RAND_2514;
  reg [31:0] _RAND_2515;
  reg [31:0] _RAND_2516;
  reg [31:0] _RAND_2517;
  reg [31:0] _RAND_2518;
  reg [31:0] _RAND_2519;
  reg [31:0] _RAND_2520;
  reg [31:0] _RAND_2521;
  reg [31:0] _RAND_2522;
  reg [31:0] _RAND_2523;
  reg [31:0] _RAND_2524;
  reg [31:0] _RAND_2525;
  reg [31:0] _RAND_2526;
  reg [31:0] _RAND_2527;
  reg [31:0] _RAND_2528;
  reg [31:0] _RAND_2529;
  reg [31:0] _RAND_2530;
  reg [31:0] _RAND_2531;
  reg [31:0] _RAND_2532;
  reg [31:0] _RAND_2533;
  reg [31:0] _RAND_2534;
  reg [31:0] _RAND_2535;
  reg [31:0] _RAND_2536;
  reg [31:0] _RAND_2537;
  reg [31:0] _RAND_2538;
  reg [31:0] _RAND_2539;
  reg [31:0] _RAND_2540;
  reg [31:0] _RAND_2541;
  reg [31:0] _RAND_2542;
  reg [31:0] _RAND_2543;
  reg [31:0] _RAND_2544;
  reg [31:0] _RAND_2545;
  reg [31:0] _RAND_2546;
  reg [31:0] _RAND_2547;
  reg [31:0] _RAND_2548;
  reg [31:0] _RAND_2549;
  reg [31:0] _RAND_2550;
  reg [31:0] _RAND_2551;
  reg [31:0] _RAND_2552;
  reg [31:0] _RAND_2553;
  reg [31:0] _RAND_2554;
  reg [31:0] _RAND_2555;
  reg [31:0] _RAND_2556;
  reg [31:0] _RAND_2557;
  reg [31:0] _RAND_2558;
  reg [31:0] _RAND_2559;
  reg [31:0] _RAND_2560;
  reg [31:0] _RAND_2561;
  reg [31:0] _RAND_2562;
  reg [31:0] _RAND_2563;
  reg [31:0] _RAND_2564;
  reg [31:0] _RAND_2565;
  reg [31:0] _RAND_2566;
  reg [31:0] _RAND_2567;
  reg [31:0] _RAND_2568;
  reg [31:0] _RAND_2569;
  reg [31:0] _RAND_2570;
  reg [31:0] _RAND_2571;
  reg [31:0] _RAND_2572;
  reg [31:0] _RAND_2573;
  reg [31:0] _RAND_2574;
  reg [31:0] _RAND_2575;
  reg [31:0] _RAND_2576;
  reg [31:0] _RAND_2577;
  reg [31:0] _RAND_2578;
  reg [31:0] _RAND_2579;
  reg [31:0] _RAND_2580;
  reg [31:0] _RAND_2581;
  reg [31:0] _RAND_2582;
  reg [31:0] _RAND_2583;
  reg [31:0] _RAND_2584;
  reg [31:0] _RAND_2585;
  reg [31:0] _RAND_2586;
  reg [31:0] _RAND_2587;
  reg [31:0] _RAND_2588;
  reg [31:0] _RAND_2589;
  reg [31:0] _RAND_2590;
  reg [31:0] _RAND_2591;
  reg [31:0] _RAND_2592;
  reg [31:0] _RAND_2593;
  reg [31:0] _RAND_2594;
  reg [31:0] _RAND_2595;
  reg [31:0] _RAND_2596;
  reg [31:0] _RAND_2597;
  reg [31:0] _RAND_2598;
  reg [31:0] _RAND_2599;
  reg [31:0] _RAND_2600;
  reg [31:0] _RAND_2601;
  reg [31:0] _RAND_2602;
  reg [31:0] _RAND_2603;
  reg [31:0] _RAND_2604;
  reg [31:0] _RAND_2605;
  reg [31:0] _RAND_2606;
  reg [31:0] _RAND_2607;
  reg [31:0] _RAND_2608;
  reg [31:0] _RAND_2609;
  reg [31:0] _RAND_2610;
  reg [31:0] _RAND_2611;
  reg [31:0] _RAND_2612;
  reg [31:0] _RAND_2613;
  reg [31:0] _RAND_2614;
  reg [31:0] _RAND_2615;
  reg [31:0] _RAND_2616;
  reg [31:0] _RAND_2617;
  reg [31:0] _RAND_2618;
  reg [31:0] _RAND_2619;
  reg [31:0] _RAND_2620;
  reg [31:0] _RAND_2621;
  reg [31:0] _RAND_2622;
  reg [31:0] _RAND_2623;
  reg [31:0] _RAND_2624;
  reg [31:0] _RAND_2625;
  reg [31:0] _RAND_2626;
  reg [31:0] _RAND_2627;
  reg [31:0] _RAND_2628;
  reg [31:0] _RAND_2629;
  reg [31:0] _RAND_2630;
  reg [31:0] _RAND_2631;
  reg [31:0] _RAND_2632;
  reg [31:0] _RAND_2633;
  reg [31:0] _RAND_2634;
  reg [31:0] _RAND_2635;
  reg [31:0] _RAND_2636;
  reg [31:0] _RAND_2637;
  reg [31:0] _RAND_2638;
  reg [31:0] _RAND_2639;
  reg [31:0] _RAND_2640;
  reg [31:0] _RAND_2641;
  reg [31:0] _RAND_2642;
  reg [31:0] _RAND_2643;
  reg [31:0] _RAND_2644;
  reg [31:0] _RAND_2645;
  reg [31:0] _RAND_2646;
  reg [31:0] _RAND_2647;
  reg [31:0] _RAND_2648;
  reg [31:0] _RAND_2649;
  reg [31:0] _RAND_2650;
  reg [31:0] _RAND_2651;
  reg [31:0] _RAND_2652;
  reg [31:0] _RAND_2653;
  reg [31:0] _RAND_2654;
  reg [31:0] _RAND_2655;
  reg [31:0] _RAND_2656;
  reg [31:0] _RAND_2657;
  reg [31:0] _RAND_2658;
  reg [31:0] _RAND_2659;
  reg [31:0] _RAND_2660;
  reg [31:0] _RAND_2661;
  reg [31:0] _RAND_2662;
  reg [31:0] _RAND_2663;
  reg [31:0] _RAND_2664;
  reg [31:0] _RAND_2665;
  reg [31:0] _RAND_2666;
  reg [31:0] _RAND_2667;
  reg [31:0] _RAND_2668;
  reg [31:0] _RAND_2669;
  reg [31:0] _RAND_2670;
  reg [31:0] _RAND_2671;
  reg [31:0] _RAND_2672;
  reg [31:0] _RAND_2673;
  reg [31:0] _RAND_2674;
  reg [31:0] _RAND_2675;
  reg [31:0] _RAND_2676;
  reg [31:0] _RAND_2677;
  reg [31:0] _RAND_2678;
  reg [31:0] _RAND_2679;
  reg [31:0] _RAND_2680;
  reg [31:0] _RAND_2681;
  reg [31:0] _RAND_2682;
  reg [31:0] _RAND_2683;
  reg [31:0] _RAND_2684;
  reg [31:0] _RAND_2685;
  reg [31:0] _RAND_2686;
  reg [31:0] _RAND_2687;
  reg [31:0] _RAND_2688;
  reg [31:0] _RAND_2689;
  reg [31:0] _RAND_2690;
  reg [31:0] _RAND_2691;
  reg [31:0] _RAND_2692;
  reg [31:0] _RAND_2693;
  reg [31:0] _RAND_2694;
  reg [31:0] _RAND_2695;
  reg [31:0] _RAND_2696;
  reg [31:0] _RAND_2697;
  reg [31:0] _RAND_2698;
  reg [31:0] _RAND_2699;
  reg [31:0] _RAND_2700;
  reg [31:0] _RAND_2701;
  reg [31:0] _RAND_2702;
  reg [31:0] _RAND_2703;
  reg [31:0] _RAND_2704;
  reg [31:0] _RAND_2705;
  reg [31:0] _RAND_2706;
  reg [31:0] _RAND_2707;
  reg [31:0] _RAND_2708;
  reg [31:0] _RAND_2709;
  reg [31:0] _RAND_2710;
  reg [31:0] _RAND_2711;
  reg [31:0] _RAND_2712;
  reg [31:0] _RAND_2713;
  reg [31:0] _RAND_2714;
  reg [31:0] _RAND_2715;
  reg [31:0] _RAND_2716;
  reg [31:0] _RAND_2717;
  reg [31:0] _RAND_2718;
  reg [31:0] _RAND_2719;
  reg [31:0] _RAND_2720;
  reg [31:0] _RAND_2721;
  reg [31:0] _RAND_2722;
  reg [31:0] _RAND_2723;
  reg [31:0] _RAND_2724;
  reg [31:0] _RAND_2725;
  reg [31:0] _RAND_2726;
  reg [31:0] _RAND_2727;
  reg [31:0] _RAND_2728;
  reg [31:0] _RAND_2729;
  reg [31:0] _RAND_2730;
  reg [31:0] _RAND_2731;
  reg [31:0] _RAND_2732;
  reg [31:0] _RAND_2733;
  reg [31:0] _RAND_2734;
  reg [31:0] _RAND_2735;
  reg [31:0] _RAND_2736;
  reg [31:0] _RAND_2737;
  reg [31:0] _RAND_2738;
  reg [31:0] _RAND_2739;
  reg [31:0] _RAND_2740;
  reg [31:0] _RAND_2741;
  reg [31:0] _RAND_2742;
  reg [31:0] _RAND_2743;
  reg [31:0] _RAND_2744;
  reg [31:0] _RAND_2745;
  reg [31:0] _RAND_2746;
  reg [31:0] _RAND_2747;
  reg [31:0] _RAND_2748;
  reg [31:0] _RAND_2749;
  reg [31:0] _RAND_2750;
  reg [31:0] _RAND_2751;
  reg [31:0] _RAND_2752;
  reg [31:0] _RAND_2753;
  reg [31:0] _RAND_2754;
  reg [31:0] _RAND_2755;
  reg [31:0] _RAND_2756;
  reg [31:0] _RAND_2757;
  reg [31:0] _RAND_2758;
  reg [31:0] _RAND_2759;
  reg [31:0] _RAND_2760;
  reg [31:0] _RAND_2761;
  reg [31:0] _RAND_2762;
  reg [31:0] _RAND_2763;
  reg [31:0] _RAND_2764;
  reg [31:0] _RAND_2765;
  reg [31:0] _RAND_2766;
  reg [31:0] _RAND_2767;
  reg [31:0] _RAND_2768;
  reg [31:0] _RAND_2769;
  reg [31:0] _RAND_2770;
  reg [31:0] _RAND_2771;
  reg [31:0] _RAND_2772;
  reg [31:0] _RAND_2773;
  reg [31:0] _RAND_2774;
  reg [31:0] _RAND_2775;
  reg [31:0] _RAND_2776;
  reg [31:0] _RAND_2777;
  reg [31:0] _RAND_2778;
  reg [31:0] _RAND_2779;
  reg [31:0] _RAND_2780;
  reg [31:0] _RAND_2781;
  reg [31:0] _RAND_2782;
  reg [31:0] _RAND_2783;
  reg [31:0] _RAND_2784;
  reg [31:0] _RAND_2785;
  reg [31:0] _RAND_2786;
  reg [31:0] _RAND_2787;
  reg [31:0] _RAND_2788;
  reg [31:0] _RAND_2789;
  reg [31:0] _RAND_2790;
  reg [31:0] _RAND_2791;
  reg [31:0] _RAND_2792;
  reg [31:0] _RAND_2793;
  reg [31:0] _RAND_2794;
  reg [31:0] _RAND_2795;
  reg [31:0] _RAND_2796;
  reg [31:0] _RAND_2797;
  reg [31:0] _RAND_2798;
  reg [31:0] _RAND_2799;
  reg [31:0] _RAND_2800;
  reg [31:0] _RAND_2801;
  reg [31:0] _RAND_2802;
  reg [31:0] _RAND_2803;
  reg [31:0] _RAND_2804;
  reg [31:0] _RAND_2805;
  reg [31:0] _RAND_2806;
  reg [31:0] _RAND_2807;
  reg [31:0] _RAND_2808;
  reg [31:0] _RAND_2809;
  reg [31:0] _RAND_2810;
  reg [31:0] _RAND_2811;
  reg [31:0] _RAND_2812;
  reg [31:0] _RAND_2813;
  reg [31:0] _RAND_2814;
  reg [31:0] _RAND_2815;
  reg [31:0] _RAND_2816;
  reg [31:0] _RAND_2817;
  reg [31:0] _RAND_2818;
  reg [31:0] _RAND_2819;
  reg [31:0] _RAND_2820;
  reg [31:0] _RAND_2821;
  reg [31:0] _RAND_2822;
  reg [31:0] _RAND_2823;
  reg [31:0] _RAND_2824;
  reg [31:0] _RAND_2825;
  reg [31:0] _RAND_2826;
  reg [31:0] _RAND_2827;
  reg [31:0] _RAND_2828;
  reg [31:0] _RAND_2829;
  reg [31:0] _RAND_2830;
  reg [31:0] _RAND_2831;
  reg [31:0] _RAND_2832;
  reg [31:0] _RAND_2833;
  reg [31:0] _RAND_2834;
  reg [31:0] _RAND_2835;
  reg [31:0] _RAND_2836;
  reg [31:0] _RAND_2837;
  reg [31:0] _RAND_2838;
  reg [31:0] _RAND_2839;
  reg [31:0] _RAND_2840;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] m_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_1_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_1_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_1_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_1_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_2_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_2_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_2_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_2_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_3_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_3_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_3_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_3_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_4_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_4_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_4_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_4_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_5_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_5_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_5_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_5_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_6_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_6_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_6_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_6_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_7_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_7_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_7_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_7_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_8_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_8_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_8_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_8_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_9_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_9_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_9_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_9_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_10_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_10_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_10_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_10_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_11_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_11_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_11_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_11_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_12_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_12_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_12_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_12_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_13_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_13_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_13_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_13_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_14_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_14_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_14_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_14_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_15_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_15_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_15_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_15_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_16_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_16_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_16_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_16_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_17_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_17_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_17_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_17_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_18_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_18_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_18_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_18_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_19_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_19_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_19_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_19_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_20_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_20_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_20_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_20_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_21_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_21_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_21_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_21_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_22_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_22_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_22_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_22_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_23_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_23_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_23_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_23_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_24_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_24_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_24_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_24_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_25_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_25_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_25_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_25_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_26_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_26_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_26_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_26_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_27_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_27_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_27_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_27_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_28_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_28_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_28_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_28_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_29_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_29_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_29_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_29_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_30_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_30_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_30_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_30_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_31_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_31_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_31_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_31_io_carry; // @[MUL.scala 81:21]
  wire [2:0] m_32_io_y_3; // @[MUL.scala 81:21]
  wire [65:0] m_32_io_x; // @[MUL.scala 81:21]
  wire [65:0] m_32_io_p; // @[MUL.scala 81:21]
  wire [1:0] m_32_io_carry; // @[MUL.scala 81:21]
  wire  m_33_io_in_0; // @[MUL.scala 124:19]
  wire  m_33_io_in_1; // @[MUL.scala 124:19]
  wire  m_33_io_out_0; // @[MUL.scala 124:19]
  wire  m_33_io_out_1; // @[MUL.scala 124:19]
  wire  m_34_io_in_0; // @[MUL.scala 124:19]
  wire  m_34_io_in_1; // @[MUL.scala 124:19]
  wire  m_34_io_out_0; // @[MUL.scala 124:19]
  wire  m_34_io_out_1; // @[MUL.scala 124:19]
  wire  m_35_io_x1; // @[MUL.scala 102:19]
  wire  m_35_io_x2; // @[MUL.scala 102:19]
  wire  m_35_io_x3; // @[MUL.scala 102:19]
  wire  m_35_io_s; // @[MUL.scala 102:19]
  wire  m_35_io_cout; // @[MUL.scala 102:19]
  wire  m_36_io_x1; // @[MUL.scala 102:19]
  wire  m_36_io_x2; // @[MUL.scala 102:19]
  wire  m_36_io_x3; // @[MUL.scala 102:19]
  wire  m_36_io_s; // @[MUL.scala 102:19]
  wire  m_36_io_cout; // @[MUL.scala 102:19]
  wire  m_37_io_x1; // @[MUL.scala 102:19]
  wire  m_37_io_x2; // @[MUL.scala 102:19]
  wire  m_37_io_x3; // @[MUL.scala 102:19]
  wire  m_37_io_s; // @[MUL.scala 102:19]
  wire  m_37_io_cout; // @[MUL.scala 102:19]
  wire  m_38_io_x1; // @[MUL.scala 102:19]
  wire  m_38_io_x2; // @[MUL.scala 102:19]
  wire  m_38_io_x3; // @[MUL.scala 102:19]
  wire  m_38_io_s; // @[MUL.scala 102:19]
  wire  m_38_io_cout; // @[MUL.scala 102:19]
  wire  m_39_io_x1; // @[MUL.scala 102:19]
  wire  m_39_io_x2; // @[MUL.scala 102:19]
  wire  m_39_io_x3; // @[MUL.scala 102:19]
  wire  m_39_io_s; // @[MUL.scala 102:19]
  wire  m_39_io_cout; // @[MUL.scala 102:19]
  wire  m_40_io_in_0; // @[MUL.scala 124:19]
  wire  m_40_io_in_1; // @[MUL.scala 124:19]
  wire  m_40_io_out_0; // @[MUL.scala 124:19]
  wire  m_40_io_out_1; // @[MUL.scala 124:19]
  wire  m_41_io_x1; // @[MUL.scala 102:19]
  wire  m_41_io_x2; // @[MUL.scala 102:19]
  wire  m_41_io_x3; // @[MUL.scala 102:19]
  wire  m_41_io_s; // @[MUL.scala 102:19]
  wire  m_41_io_cout; // @[MUL.scala 102:19]
  wire  m_42_io_in_0; // @[MUL.scala 124:19]
  wire  m_42_io_in_1; // @[MUL.scala 124:19]
  wire  m_42_io_out_0; // @[MUL.scala 124:19]
  wire  m_42_io_out_1; // @[MUL.scala 124:19]
  wire  m_43_io_x1; // @[MUL.scala 102:19]
  wire  m_43_io_x2; // @[MUL.scala 102:19]
  wire  m_43_io_x3; // @[MUL.scala 102:19]
  wire  m_43_io_s; // @[MUL.scala 102:19]
  wire  m_43_io_cout; // @[MUL.scala 102:19]
  wire  m_44_io_x1; // @[MUL.scala 102:19]
  wire  m_44_io_x2; // @[MUL.scala 102:19]
  wire  m_44_io_x3; // @[MUL.scala 102:19]
  wire  m_44_io_s; // @[MUL.scala 102:19]
  wire  m_44_io_cout; // @[MUL.scala 102:19]
  wire  m_45_io_x1; // @[MUL.scala 102:19]
  wire  m_45_io_x2; // @[MUL.scala 102:19]
  wire  m_45_io_x3; // @[MUL.scala 102:19]
  wire  m_45_io_s; // @[MUL.scala 102:19]
  wire  m_45_io_cout; // @[MUL.scala 102:19]
  wire  m_46_io_x1; // @[MUL.scala 102:19]
  wire  m_46_io_x2; // @[MUL.scala 102:19]
  wire  m_46_io_x3; // @[MUL.scala 102:19]
  wire  m_46_io_s; // @[MUL.scala 102:19]
  wire  m_46_io_cout; // @[MUL.scala 102:19]
  wire  m_47_io_x1; // @[MUL.scala 102:19]
  wire  m_47_io_x2; // @[MUL.scala 102:19]
  wire  m_47_io_x3; // @[MUL.scala 102:19]
  wire  m_47_io_s; // @[MUL.scala 102:19]
  wire  m_47_io_cout; // @[MUL.scala 102:19]
  wire  m_48_io_x1; // @[MUL.scala 102:19]
  wire  m_48_io_x2; // @[MUL.scala 102:19]
  wire  m_48_io_x3; // @[MUL.scala 102:19]
  wire  m_48_io_s; // @[MUL.scala 102:19]
  wire  m_48_io_cout; // @[MUL.scala 102:19]
  wire  m_49_io_x1; // @[MUL.scala 102:19]
  wire  m_49_io_x2; // @[MUL.scala 102:19]
  wire  m_49_io_x3; // @[MUL.scala 102:19]
  wire  m_49_io_s; // @[MUL.scala 102:19]
  wire  m_49_io_cout; // @[MUL.scala 102:19]
  wire  m_50_io_x1; // @[MUL.scala 102:19]
  wire  m_50_io_x2; // @[MUL.scala 102:19]
  wire  m_50_io_x3; // @[MUL.scala 102:19]
  wire  m_50_io_s; // @[MUL.scala 102:19]
  wire  m_50_io_cout; // @[MUL.scala 102:19]
  wire  m_51_io_x1; // @[MUL.scala 102:19]
  wire  m_51_io_x2; // @[MUL.scala 102:19]
  wire  m_51_io_x3; // @[MUL.scala 102:19]
  wire  m_51_io_s; // @[MUL.scala 102:19]
  wire  m_51_io_cout; // @[MUL.scala 102:19]
  wire  m_52_io_x1; // @[MUL.scala 102:19]
  wire  m_52_io_x2; // @[MUL.scala 102:19]
  wire  m_52_io_x3; // @[MUL.scala 102:19]
  wire  m_52_io_s; // @[MUL.scala 102:19]
  wire  m_52_io_cout; // @[MUL.scala 102:19]
  wire  m_53_io_in_0; // @[MUL.scala 124:19]
  wire  m_53_io_in_1; // @[MUL.scala 124:19]
  wire  m_53_io_out_0; // @[MUL.scala 124:19]
  wire  m_53_io_out_1; // @[MUL.scala 124:19]
  wire  m_54_io_x1; // @[MUL.scala 102:19]
  wire  m_54_io_x2; // @[MUL.scala 102:19]
  wire  m_54_io_x3; // @[MUL.scala 102:19]
  wire  m_54_io_s; // @[MUL.scala 102:19]
  wire  m_54_io_cout; // @[MUL.scala 102:19]
  wire  m_55_io_x1; // @[MUL.scala 102:19]
  wire  m_55_io_x2; // @[MUL.scala 102:19]
  wire  m_55_io_x3; // @[MUL.scala 102:19]
  wire  m_55_io_s; // @[MUL.scala 102:19]
  wire  m_55_io_cout; // @[MUL.scala 102:19]
  wire  m_56_io_in_0; // @[MUL.scala 124:19]
  wire  m_56_io_in_1; // @[MUL.scala 124:19]
  wire  m_56_io_out_0; // @[MUL.scala 124:19]
  wire  m_56_io_out_1; // @[MUL.scala 124:19]
  wire  m_57_io_x1; // @[MUL.scala 102:19]
  wire  m_57_io_x2; // @[MUL.scala 102:19]
  wire  m_57_io_x3; // @[MUL.scala 102:19]
  wire  m_57_io_s; // @[MUL.scala 102:19]
  wire  m_57_io_cout; // @[MUL.scala 102:19]
  wire  m_58_io_x1; // @[MUL.scala 102:19]
  wire  m_58_io_x2; // @[MUL.scala 102:19]
  wire  m_58_io_x3; // @[MUL.scala 102:19]
  wire  m_58_io_s; // @[MUL.scala 102:19]
  wire  m_58_io_cout; // @[MUL.scala 102:19]
  wire  m_59_io_x1; // @[MUL.scala 102:19]
  wire  m_59_io_x2; // @[MUL.scala 102:19]
  wire  m_59_io_x3; // @[MUL.scala 102:19]
  wire  m_59_io_s; // @[MUL.scala 102:19]
  wire  m_59_io_cout; // @[MUL.scala 102:19]
  wire  m_60_io_x1; // @[MUL.scala 102:19]
  wire  m_60_io_x2; // @[MUL.scala 102:19]
  wire  m_60_io_x3; // @[MUL.scala 102:19]
  wire  m_60_io_s; // @[MUL.scala 102:19]
  wire  m_60_io_cout; // @[MUL.scala 102:19]
  wire  m_61_io_x1; // @[MUL.scala 102:19]
  wire  m_61_io_x2; // @[MUL.scala 102:19]
  wire  m_61_io_x3; // @[MUL.scala 102:19]
  wire  m_61_io_s; // @[MUL.scala 102:19]
  wire  m_61_io_cout; // @[MUL.scala 102:19]
  wire  m_62_io_x1; // @[MUL.scala 102:19]
  wire  m_62_io_x2; // @[MUL.scala 102:19]
  wire  m_62_io_x3; // @[MUL.scala 102:19]
  wire  m_62_io_s; // @[MUL.scala 102:19]
  wire  m_62_io_cout; // @[MUL.scala 102:19]
  wire  m_63_io_x1; // @[MUL.scala 102:19]
  wire  m_63_io_x2; // @[MUL.scala 102:19]
  wire  m_63_io_x3; // @[MUL.scala 102:19]
  wire  m_63_io_s; // @[MUL.scala 102:19]
  wire  m_63_io_cout; // @[MUL.scala 102:19]
  wire  m_64_io_x1; // @[MUL.scala 102:19]
  wire  m_64_io_x2; // @[MUL.scala 102:19]
  wire  m_64_io_x3; // @[MUL.scala 102:19]
  wire  m_64_io_s; // @[MUL.scala 102:19]
  wire  m_64_io_cout; // @[MUL.scala 102:19]
  wire  m_65_io_x1; // @[MUL.scala 102:19]
  wire  m_65_io_x2; // @[MUL.scala 102:19]
  wire  m_65_io_x3; // @[MUL.scala 102:19]
  wire  m_65_io_s; // @[MUL.scala 102:19]
  wire  m_65_io_cout; // @[MUL.scala 102:19]
  wire  m_66_io_x1; // @[MUL.scala 102:19]
  wire  m_66_io_x2; // @[MUL.scala 102:19]
  wire  m_66_io_x3; // @[MUL.scala 102:19]
  wire  m_66_io_s; // @[MUL.scala 102:19]
  wire  m_66_io_cout; // @[MUL.scala 102:19]
  wire  m_67_io_x1; // @[MUL.scala 102:19]
  wire  m_67_io_x2; // @[MUL.scala 102:19]
  wire  m_67_io_x3; // @[MUL.scala 102:19]
  wire  m_67_io_s; // @[MUL.scala 102:19]
  wire  m_67_io_cout; // @[MUL.scala 102:19]
  wire  m_68_io_x1; // @[MUL.scala 102:19]
  wire  m_68_io_x2; // @[MUL.scala 102:19]
  wire  m_68_io_x3; // @[MUL.scala 102:19]
  wire  m_68_io_s; // @[MUL.scala 102:19]
  wire  m_68_io_cout; // @[MUL.scala 102:19]
  wire  m_69_io_x1; // @[MUL.scala 102:19]
  wire  m_69_io_x2; // @[MUL.scala 102:19]
  wire  m_69_io_x3; // @[MUL.scala 102:19]
  wire  m_69_io_s; // @[MUL.scala 102:19]
  wire  m_69_io_cout; // @[MUL.scala 102:19]
  wire  m_70_io_x1; // @[MUL.scala 102:19]
  wire  m_70_io_x2; // @[MUL.scala 102:19]
  wire  m_70_io_x3; // @[MUL.scala 102:19]
  wire  m_70_io_s; // @[MUL.scala 102:19]
  wire  m_70_io_cout; // @[MUL.scala 102:19]
  wire  m_71_io_x1; // @[MUL.scala 102:19]
  wire  m_71_io_x2; // @[MUL.scala 102:19]
  wire  m_71_io_x3; // @[MUL.scala 102:19]
  wire  m_71_io_s; // @[MUL.scala 102:19]
  wire  m_71_io_cout; // @[MUL.scala 102:19]
  wire  m_72_io_in_0; // @[MUL.scala 124:19]
  wire  m_72_io_in_1; // @[MUL.scala 124:19]
  wire  m_72_io_out_0; // @[MUL.scala 124:19]
  wire  m_72_io_out_1; // @[MUL.scala 124:19]
  wire  m_73_io_x1; // @[MUL.scala 102:19]
  wire  m_73_io_x2; // @[MUL.scala 102:19]
  wire  m_73_io_x3; // @[MUL.scala 102:19]
  wire  m_73_io_s; // @[MUL.scala 102:19]
  wire  m_73_io_cout; // @[MUL.scala 102:19]
  wire  m_74_io_x1; // @[MUL.scala 102:19]
  wire  m_74_io_x2; // @[MUL.scala 102:19]
  wire  m_74_io_x3; // @[MUL.scala 102:19]
  wire  m_74_io_s; // @[MUL.scala 102:19]
  wire  m_74_io_cout; // @[MUL.scala 102:19]
  wire  m_75_io_x1; // @[MUL.scala 102:19]
  wire  m_75_io_x2; // @[MUL.scala 102:19]
  wire  m_75_io_x3; // @[MUL.scala 102:19]
  wire  m_75_io_s; // @[MUL.scala 102:19]
  wire  m_75_io_cout; // @[MUL.scala 102:19]
  wire  m_76_io_in_0; // @[MUL.scala 124:19]
  wire  m_76_io_in_1; // @[MUL.scala 124:19]
  wire  m_76_io_out_0; // @[MUL.scala 124:19]
  wire  m_76_io_out_1; // @[MUL.scala 124:19]
  wire  m_77_io_x1; // @[MUL.scala 102:19]
  wire  m_77_io_x2; // @[MUL.scala 102:19]
  wire  m_77_io_x3; // @[MUL.scala 102:19]
  wire  m_77_io_s; // @[MUL.scala 102:19]
  wire  m_77_io_cout; // @[MUL.scala 102:19]
  wire  m_78_io_x1; // @[MUL.scala 102:19]
  wire  m_78_io_x2; // @[MUL.scala 102:19]
  wire  m_78_io_x3; // @[MUL.scala 102:19]
  wire  m_78_io_s; // @[MUL.scala 102:19]
  wire  m_78_io_cout; // @[MUL.scala 102:19]
  wire  m_79_io_x1; // @[MUL.scala 102:19]
  wire  m_79_io_x2; // @[MUL.scala 102:19]
  wire  m_79_io_x3; // @[MUL.scala 102:19]
  wire  m_79_io_s; // @[MUL.scala 102:19]
  wire  m_79_io_cout; // @[MUL.scala 102:19]
  wire  m_80_io_x1; // @[MUL.scala 102:19]
  wire  m_80_io_x2; // @[MUL.scala 102:19]
  wire  m_80_io_x3; // @[MUL.scala 102:19]
  wire  m_80_io_s; // @[MUL.scala 102:19]
  wire  m_80_io_cout; // @[MUL.scala 102:19]
  wire  m_81_io_x1; // @[MUL.scala 102:19]
  wire  m_81_io_x2; // @[MUL.scala 102:19]
  wire  m_81_io_x3; // @[MUL.scala 102:19]
  wire  m_81_io_s; // @[MUL.scala 102:19]
  wire  m_81_io_cout; // @[MUL.scala 102:19]
  wire  m_82_io_x1; // @[MUL.scala 102:19]
  wire  m_82_io_x2; // @[MUL.scala 102:19]
  wire  m_82_io_x3; // @[MUL.scala 102:19]
  wire  m_82_io_s; // @[MUL.scala 102:19]
  wire  m_82_io_cout; // @[MUL.scala 102:19]
  wire  m_83_io_x1; // @[MUL.scala 102:19]
  wire  m_83_io_x2; // @[MUL.scala 102:19]
  wire  m_83_io_x3; // @[MUL.scala 102:19]
  wire  m_83_io_s; // @[MUL.scala 102:19]
  wire  m_83_io_cout; // @[MUL.scala 102:19]
  wire  m_84_io_x1; // @[MUL.scala 102:19]
  wire  m_84_io_x2; // @[MUL.scala 102:19]
  wire  m_84_io_x3; // @[MUL.scala 102:19]
  wire  m_84_io_s; // @[MUL.scala 102:19]
  wire  m_84_io_cout; // @[MUL.scala 102:19]
  wire  m_85_io_x1; // @[MUL.scala 102:19]
  wire  m_85_io_x2; // @[MUL.scala 102:19]
  wire  m_85_io_x3; // @[MUL.scala 102:19]
  wire  m_85_io_s; // @[MUL.scala 102:19]
  wire  m_85_io_cout; // @[MUL.scala 102:19]
  wire  m_86_io_x1; // @[MUL.scala 102:19]
  wire  m_86_io_x2; // @[MUL.scala 102:19]
  wire  m_86_io_x3; // @[MUL.scala 102:19]
  wire  m_86_io_s; // @[MUL.scala 102:19]
  wire  m_86_io_cout; // @[MUL.scala 102:19]
  wire  m_87_io_x1; // @[MUL.scala 102:19]
  wire  m_87_io_x2; // @[MUL.scala 102:19]
  wire  m_87_io_x3; // @[MUL.scala 102:19]
  wire  m_87_io_s; // @[MUL.scala 102:19]
  wire  m_87_io_cout; // @[MUL.scala 102:19]
  wire  m_88_io_x1; // @[MUL.scala 102:19]
  wire  m_88_io_x2; // @[MUL.scala 102:19]
  wire  m_88_io_x3; // @[MUL.scala 102:19]
  wire  m_88_io_s; // @[MUL.scala 102:19]
  wire  m_88_io_cout; // @[MUL.scala 102:19]
  wire  m_89_io_x1; // @[MUL.scala 102:19]
  wire  m_89_io_x2; // @[MUL.scala 102:19]
  wire  m_89_io_x3; // @[MUL.scala 102:19]
  wire  m_89_io_s; // @[MUL.scala 102:19]
  wire  m_89_io_cout; // @[MUL.scala 102:19]
  wire  m_90_io_x1; // @[MUL.scala 102:19]
  wire  m_90_io_x2; // @[MUL.scala 102:19]
  wire  m_90_io_x3; // @[MUL.scala 102:19]
  wire  m_90_io_s; // @[MUL.scala 102:19]
  wire  m_90_io_cout; // @[MUL.scala 102:19]
  wire  m_91_io_x1; // @[MUL.scala 102:19]
  wire  m_91_io_x2; // @[MUL.scala 102:19]
  wire  m_91_io_x3; // @[MUL.scala 102:19]
  wire  m_91_io_s; // @[MUL.scala 102:19]
  wire  m_91_io_cout; // @[MUL.scala 102:19]
  wire  m_92_io_x1; // @[MUL.scala 102:19]
  wire  m_92_io_x2; // @[MUL.scala 102:19]
  wire  m_92_io_x3; // @[MUL.scala 102:19]
  wire  m_92_io_s; // @[MUL.scala 102:19]
  wire  m_92_io_cout; // @[MUL.scala 102:19]
  wire  m_93_io_x1; // @[MUL.scala 102:19]
  wire  m_93_io_x2; // @[MUL.scala 102:19]
  wire  m_93_io_x3; // @[MUL.scala 102:19]
  wire  m_93_io_s; // @[MUL.scala 102:19]
  wire  m_93_io_cout; // @[MUL.scala 102:19]
  wire  m_94_io_x1; // @[MUL.scala 102:19]
  wire  m_94_io_x2; // @[MUL.scala 102:19]
  wire  m_94_io_x3; // @[MUL.scala 102:19]
  wire  m_94_io_s; // @[MUL.scala 102:19]
  wire  m_94_io_cout; // @[MUL.scala 102:19]
  wire  m_95_io_x1; // @[MUL.scala 102:19]
  wire  m_95_io_x2; // @[MUL.scala 102:19]
  wire  m_95_io_x3; // @[MUL.scala 102:19]
  wire  m_95_io_s; // @[MUL.scala 102:19]
  wire  m_95_io_cout; // @[MUL.scala 102:19]
  wire  m_96_io_x1; // @[MUL.scala 102:19]
  wire  m_96_io_x2; // @[MUL.scala 102:19]
  wire  m_96_io_x3; // @[MUL.scala 102:19]
  wire  m_96_io_s; // @[MUL.scala 102:19]
  wire  m_96_io_cout; // @[MUL.scala 102:19]
  wire  m_97_io_in_0; // @[MUL.scala 124:19]
  wire  m_97_io_in_1; // @[MUL.scala 124:19]
  wire  m_97_io_out_0; // @[MUL.scala 124:19]
  wire  m_97_io_out_1; // @[MUL.scala 124:19]
  wire  m_98_io_x1; // @[MUL.scala 102:19]
  wire  m_98_io_x2; // @[MUL.scala 102:19]
  wire  m_98_io_x3; // @[MUL.scala 102:19]
  wire  m_98_io_s; // @[MUL.scala 102:19]
  wire  m_98_io_cout; // @[MUL.scala 102:19]
  wire  m_99_io_x1; // @[MUL.scala 102:19]
  wire  m_99_io_x2; // @[MUL.scala 102:19]
  wire  m_99_io_x3; // @[MUL.scala 102:19]
  wire  m_99_io_s; // @[MUL.scala 102:19]
  wire  m_99_io_cout; // @[MUL.scala 102:19]
  wire  m_100_io_x1; // @[MUL.scala 102:19]
  wire  m_100_io_x2; // @[MUL.scala 102:19]
  wire  m_100_io_x3; // @[MUL.scala 102:19]
  wire  m_100_io_s; // @[MUL.scala 102:19]
  wire  m_100_io_cout; // @[MUL.scala 102:19]
  wire  m_101_io_x1; // @[MUL.scala 102:19]
  wire  m_101_io_x2; // @[MUL.scala 102:19]
  wire  m_101_io_x3; // @[MUL.scala 102:19]
  wire  m_101_io_s; // @[MUL.scala 102:19]
  wire  m_101_io_cout; // @[MUL.scala 102:19]
  wire  m_102_io_in_0; // @[MUL.scala 124:19]
  wire  m_102_io_in_1; // @[MUL.scala 124:19]
  wire  m_102_io_out_0; // @[MUL.scala 124:19]
  wire  m_102_io_out_1; // @[MUL.scala 124:19]
  wire  m_103_io_x1; // @[MUL.scala 102:19]
  wire  m_103_io_x2; // @[MUL.scala 102:19]
  wire  m_103_io_x3; // @[MUL.scala 102:19]
  wire  m_103_io_s; // @[MUL.scala 102:19]
  wire  m_103_io_cout; // @[MUL.scala 102:19]
  wire  m_104_io_x1; // @[MUL.scala 102:19]
  wire  m_104_io_x2; // @[MUL.scala 102:19]
  wire  m_104_io_x3; // @[MUL.scala 102:19]
  wire  m_104_io_s; // @[MUL.scala 102:19]
  wire  m_104_io_cout; // @[MUL.scala 102:19]
  wire  m_105_io_x1; // @[MUL.scala 102:19]
  wire  m_105_io_x2; // @[MUL.scala 102:19]
  wire  m_105_io_x3; // @[MUL.scala 102:19]
  wire  m_105_io_s; // @[MUL.scala 102:19]
  wire  m_105_io_cout; // @[MUL.scala 102:19]
  wire  m_106_io_x1; // @[MUL.scala 102:19]
  wire  m_106_io_x2; // @[MUL.scala 102:19]
  wire  m_106_io_x3; // @[MUL.scala 102:19]
  wire  m_106_io_s; // @[MUL.scala 102:19]
  wire  m_106_io_cout; // @[MUL.scala 102:19]
  wire  m_107_io_x1; // @[MUL.scala 102:19]
  wire  m_107_io_x2; // @[MUL.scala 102:19]
  wire  m_107_io_x3; // @[MUL.scala 102:19]
  wire  m_107_io_s; // @[MUL.scala 102:19]
  wire  m_107_io_cout; // @[MUL.scala 102:19]
  wire  m_108_io_x1; // @[MUL.scala 102:19]
  wire  m_108_io_x2; // @[MUL.scala 102:19]
  wire  m_108_io_x3; // @[MUL.scala 102:19]
  wire  m_108_io_s; // @[MUL.scala 102:19]
  wire  m_108_io_cout; // @[MUL.scala 102:19]
  wire  m_109_io_x1; // @[MUL.scala 102:19]
  wire  m_109_io_x2; // @[MUL.scala 102:19]
  wire  m_109_io_x3; // @[MUL.scala 102:19]
  wire  m_109_io_s; // @[MUL.scala 102:19]
  wire  m_109_io_cout; // @[MUL.scala 102:19]
  wire  m_110_io_x1; // @[MUL.scala 102:19]
  wire  m_110_io_x2; // @[MUL.scala 102:19]
  wire  m_110_io_x3; // @[MUL.scala 102:19]
  wire  m_110_io_s; // @[MUL.scala 102:19]
  wire  m_110_io_cout; // @[MUL.scala 102:19]
  wire  m_111_io_x1; // @[MUL.scala 102:19]
  wire  m_111_io_x2; // @[MUL.scala 102:19]
  wire  m_111_io_x3; // @[MUL.scala 102:19]
  wire  m_111_io_s; // @[MUL.scala 102:19]
  wire  m_111_io_cout; // @[MUL.scala 102:19]
  wire  m_112_io_x1; // @[MUL.scala 102:19]
  wire  m_112_io_x2; // @[MUL.scala 102:19]
  wire  m_112_io_x3; // @[MUL.scala 102:19]
  wire  m_112_io_s; // @[MUL.scala 102:19]
  wire  m_112_io_cout; // @[MUL.scala 102:19]
  wire  m_113_io_x1; // @[MUL.scala 102:19]
  wire  m_113_io_x2; // @[MUL.scala 102:19]
  wire  m_113_io_x3; // @[MUL.scala 102:19]
  wire  m_113_io_s; // @[MUL.scala 102:19]
  wire  m_113_io_cout; // @[MUL.scala 102:19]
  wire  m_114_io_x1; // @[MUL.scala 102:19]
  wire  m_114_io_x2; // @[MUL.scala 102:19]
  wire  m_114_io_x3; // @[MUL.scala 102:19]
  wire  m_114_io_s; // @[MUL.scala 102:19]
  wire  m_114_io_cout; // @[MUL.scala 102:19]
  wire  m_115_io_x1; // @[MUL.scala 102:19]
  wire  m_115_io_x2; // @[MUL.scala 102:19]
  wire  m_115_io_x3; // @[MUL.scala 102:19]
  wire  m_115_io_s; // @[MUL.scala 102:19]
  wire  m_115_io_cout; // @[MUL.scala 102:19]
  wire  m_116_io_x1; // @[MUL.scala 102:19]
  wire  m_116_io_x2; // @[MUL.scala 102:19]
  wire  m_116_io_x3; // @[MUL.scala 102:19]
  wire  m_116_io_s; // @[MUL.scala 102:19]
  wire  m_116_io_cout; // @[MUL.scala 102:19]
  wire  m_117_io_x1; // @[MUL.scala 102:19]
  wire  m_117_io_x2; // @[MUL.scala 102:19]
  wire  m_117_io_x3; // @[MUL.scala 102:19]
  wire  m_117_io_s; // @[MUL.scala 102:19]
  wire  m_117_io_cout; // @[MUL.scala 102:19]
  wire  m_118_io_x1; // @[MUL.scala 102:19]
  wire  m_118_io_x2; // @[MUL.scala 102:19]
  wire  m_118_io_x3; // @[MUL.scala 102:19]
  wire  m_118_io_s; // @[MUL.scala 102:19]
  wire  m_118_io_cout; // @[MUL.scala 102:19]
  wire  m_119_io_x1; // @[MUL.scala 102:19]
  wire  m_119_io_x2; // @[MUL.scala 102:19]
  wire  m_119_io_x3; // @[MUL.scala 102:19]
  wire  m_119_io_s; // @[MUL.scala 102:19]
  wire  m_119_io_cout; // @[MUL.scala 102:19]
  wire  m_120_io_x1; // @[MUL.scala 102:19]
  wire  m_120_io_x2; // @[MUL.scala 102:19]
  wire  m_120_io_x3; // @[MUL.scala 102:19]
  wire  m_120_io_s; // @[MUL.scala 102:19]
  wire  m_120_io_cout; // @[MUL.scala 102:19]
  wire  m_121_io_x1; // @[MUL.scala 102:19]
  wire  m_121_io_x2; // @[MUL.scala 102:19]
  wire  m_121_io_x3; // @[MUL.scala 102:19]
  wire  m_121_io_s; // @[MUL.scala 102:19]
  wire  m_121_io_cout; // @[MUL.scala 102:19]
  wire  m_122_io_x1; // @[MUL.scala 102:19]
  wire  m_122_io_x2; // @[MUL.scala 102:19]
  wire  m_122_io_x3; // @[MUL.scala 102:19]
  wire  m_122_io_s; // @[MUL.scala 102:19]
  wire  m_122_io_cout; // @[MUL.scala 102:19]
  wire  m_123_io_x1; // @[MUL.scala 102:19]
  wire  m_123_io_x2; // @[MUL.scala 102:19]
  wire  m_123_io_x3; // @[MUL.scala 102:19]
  wire  m_123_io_s; // @[MUL.scala 102:19]
  wire  m_123_io_cout; // @[MUL.scala 102:19]
  wire  m_124_io_x1; // @[MUL.scala 102:19]
  wire  m_124_io_x2; // @[MUL.scala 102:19]
  wire  m_124_io_x3; // @[MUL.scala 102:19]
  wire  m_124_io_s; // @[MUL.scala 102:19]
  wire  m_124_io_cout; // @[MUL.scala 102:19]
  wire  m_125_io_x1; // @[MUL.scala 102:19]
  wire  m_125_io_x2; // @[MUL.scala 102:19]
  wire  m_125_io_x3; // @[MUL.scala 102:19]
  wire  m_125_io_s; // @[MUL.scala 102:19]
  wire  m_125_io_cout; // @[MUL.scala 102:19]
  wire  m_126_io_x1; // @[MUL.scala 102:19]
  wire  m_126_io_x2; // @[MUL.scala 102:19]
  wire  m_126_io_x3; // @[MUL.scala 102:19]
  wire  m_126_io_s; // @[MUL.scala 102:19]
  wire  m_126_io_cout; // @[MUL.scala 102:19]
  wire  m_127_io_x1; // @[MUL.scala 102:19]
  wire  m_127_io_x2; // @[MUL.scala 102:19]
  wire  m_127_io_x3; // @[MUL.scala 102:19]
  wire  m_127_io_s; // @[MUL.scala 102:19]
  wire  m_127_io_cout; // @[MUL.scala 102:19]
  wire  m_128_io_in_0; // @[MUL.scala 124:19]
  wire  m_128_io_in_1; // @[MUL.scala 124:19]
  wire  m_128_io_out_0; // @[MUL.scala 124:19]
  wire  m_128_io_out_1; // @[MUL.scala 124:19]
  wire  m_129_io_x1; // @[MUL.scala 102:19]
  wire  m_129_io_x2; // @[MUL.scala 102:19]
  wire  m_129_io_x3; // @[MUL.scala 102:19]
  wire  m_129_io_s; // @[MUL.scala 102:19]
  wire  m_129_io_cout; // @[MUL.scala 102:19]
  wire  m_130_io_x1; // @[MUL.scala 102:19]
  wire  m_130_io_x2; // @[MUL.scala 102:19]
  wire  m_130_io_x3; // @[MUL.scala 102:19]
  wire  m_130_io_s; // @[MUL.scala 102:19]
  wire  m_130_io_cout; // @[MUL.scala 102:19]
  wire  m_131_io_x1; // @[MUL.scala 102:19]
  wire  m_131_io_x2; // @[MUL.scala 102:19]
  wire  m_131_io_x3; // @[MUL.scala 102:19]
  wire  m_131_io_s; // @[MUL.scala 102:19]
  wire  m_131_io_cout; // @[MUL.scala 102:19]
  wire  m_132_io_x1; // @[MUL.scala 102:19]
  wire  m_132_io_x2; // @[MUL.scala 102:19]
  wire  m_132_io_x3; // @[MUL.scala 102:19]
  wire  m_132_io_s; // @[MUL.scala 102:19]
  wire  m_132_io_cout; // @[MUL.scala 102:19]
  wire  m_133_io_x1; // @[MUL.scala 102:19]
  wire  m_133_io_x2; // @[MUL.scala 102:19]
  wire  m_133_io_x3; // @[MUL.scala 102:19]
  wire  m_133_io_s; // @[MUL.scala 102:19]
  wire  m_133_io_cout; // @[MUL.scala 102:19]
  wire  m_134_io_in_0; // @[MUL.scala 124:19]
  wire  m_134_io_in_1; // @[MUL.scala 124:19]
  wire  m_134_io_out_0; // @[MUL.scala 124:19]
  wire  m_134_io_out_1; // @[MUL.scala 124:19]
  wire  m_135_io_x1; // @[MUL.scala 102:19]
  wire  m_135_io_x2; // @[MUL.scala 102:19]
  wire  m_135_io_x3; // @[MUL.scala 102:19]
  wire  m_135_io_s; // @[MUL.scala 102:19]
  wire  m_135_io_cout; // @[MUL.scala 102:19]
  wire  m_136_io_x1; // @[MUL.scala 102:19]
  wire  m_136_io_x2; // @[MUL.scala 102:19]
  wire  m_136_io_x3; // @[MUL.scala 102:19]
  wire  m_136_io_s; // @[MUL.scala 102:19]
  wire  m_136_io_cout; // @[MUL.scala 102:19]
  wire  m_137_io_x1; // @[MUL.scala 102:19]
  wire  m_137_io_x2; // @[MUL.scala 102:19]
  wire  m_137_io_x3; // @[MUL.scala 102:19]
  wire  m_137_io_s; // @[MUL.scala 102:19]
  wire  m_137_io_cout; // @[MUL.scala 102:19]
  wire  m_138_io_x1; // @[MUL.scala 102:19]
  wire  m_138_io_x2; // @[MUL.scala 102:19]
  wire  m_138_io_x3; // @[MUL.scala 102:19]
  wire  m_138_io_s; // @[MUL.scala 102:19]
  wire  m_138_io_cout; // @[MUL.scala 102:19]
  wire  m_139_io_x1; // @[MUL.scala 102:19]
  wire  m_139_io_x2; // @[MUL.scala 102:19]
  wire  m_139_io_x3; // @[MUL.scala 102:19]
  wire  m_139_io_s; // @[MUL.scala 102:19]
  wire  m_139_io_cout; // @[MUL.scala 102:19]
  wire  m_140_io_x1; // @[MUL.scala 102:19]
  wire  m_140_io_x2; // @[MUL.scala 102:19]
  wire  m_140_io_x3; // @[MUL.scala 102:19]
  wire  m_140_io_s; // @[MUL.scala 102:19]
  wire  m_140_io_cout; // @[MUL.scala 102:19]
  wire  m_141_io_x1; // @[MUL.scala 102:19]
  wire  m_141_io_x2; // @[MUL.scala 102:19]
  wire  m_141_io_x3; // @[MUL.scala 102:19]
  wire  m_141_io_s; // @[MUL.scala 102:19]
  wire  m_141_io_cout; // @[MUL.scala 102:19]
  wire  m_142_io_x1; // @[MUL.scala 102:19]
  wire  m_142_io_x2; // @[MUL.scala 102:19]
  wire  m_142_io_x3; // @[MUL.scala 102:19]
  wire  m_142_io_s; // @[MUL.scala 102:19]
  wire  m_142_io_cout; // @[MUL.scala 102:19]
  wire  m_143_io_x1; // @[MUL.scala 102:19]
  wire  m_143_io_x2; // @[MUL.scala 102:19]
  wire  m_143_io_x3; // @[MUL.scala 102:19]
  wire  m_143_io_s; // @[MUL.scala 102:19]
  wire  m_143_io_cout; // @[MUL.scala 102:19]
  wire  m_144_io_x1; // @[MUL.scala 102:19]
  wire  m_144_io_x2; // @[MUL.scala 102:19]
  wire  m_144_io_x3; // @[MUL.scala 102:19]
  wire  m_144_io_s; // @[MUL.scala 102:19]
  wire  m_144_io_cout; // @[MUL.scala 102:19]
  wire  m_145_io_x1; // @[MUL.scala 102:19]
  wire  m_145_io_x2; // @[MUL.scala 102:19]
  wire  m_145_io_x3; // @[MUL.scala 102:19]
  wire  m_145_io_s; // @[MUL.scala 102:19]
  wire  m_145_io_cout; // @[MUL.scala 102:19]
  wire  m_146_io_x1; // @[MUL.scala 102:19]
  wire  m_146_io_x2; // @[MUL.scala 102:19]
  wire  m_146_io_x3; // @[MUL.scala 102:19]
  wire  m_146_io_s; // @[MUL.scala 102:19]
  wire  m_146_io_cout; // @[MUL.scala 102:19]
  wire  m_147_io_x1; // @[MUL.scala 102:19]
  wire  m_147_io_x2; // @[MUL.scala 102:19]
  wire  m_147_io_x3; // @[MUL.scala 102:19]
  wire  m_147_io_s; // @[MUL.scala 102:19]
  wire  m_147_io_cout; // @[MUL.scala 102:19]
  wire  m_148_io_x1; // @[MUL.scala 102:19]
  wire  m_148_io_x2; // @[MUL.scala 102:19]
  wire  m_148_io_x3; // @[MUL.scala 102:19]
  wire  m_148_io_s; // @[MUL.scala 102:19]
  wire  m_148_io_cout; // @[MUL.scala 102:19]
  wire  m_149_io_x1; // @[MUL.scala 102:19]
  wire  m_149_io_x2; // @[MUL.scala 102:19]
  wire  m_149_io_x3; // @[MUL.scala 102:19]
  wire  m_149_io_s; // @[MUL.scala 102:19]
  wire  m_149_io_cout; // @[MUL.scala 102:19]
  wire  m_150_io_x1; // @[MUL.scala 102:19]
  wire  m_150_io_x2; // @[MUL.scala 102:19]
  wire  m_150_io_x3; // @[MUL.scala 102:19]
  wire  m_150_io_s; // @[MUL.scala 102:19]
  wire  m_150_io_cout; // @[MUL.scala 102:19]
  wire  m_151_io_x1; // @[MUL.scala 102:19]
  wire  m_151_io_x2; // @[MUL.scala 102:19]
  wire  m_151_io_x3; // @[MUL.scala 102:19]
  wire  m_151_io_s; // @[MUL.scala 102:19]
  wire  m_151_io_cout; // @[MUL.scala 102:19]
  wire  m_152_io_x1; // @[MUL.scala 102:19]
  wire  m_152_io_x2; // @[MUL.scala 102:19]
  wire  m_152_io_x3; // @[MUL.scala 102:19]
  wire  m_152_io_s; // @[MUL.scala 102:19]
  wire  m_152_io_cout; // @[MUL.scala 102:19]
  wire  m_153_io_x1; // @[MUL.scala 102:19]
  wire  m_153_io_x2; // @[MUL.scala 102:19]
  wire  m_153_io_x3; // @[MUL.scala 102:19]
  wire  m_153_io_s; // @[MUL.scala 102:19]
  wire  m_153_io_cout; // @[MUL.scala 102:19]
  wire  m_154_io_x1; // @[MUL.scala 102:19]
  wire  m_154_io_x2; // @[MUL.scala 102:19]
  wire  m_154_io_x3; // @[MUL.scala 102:19]
  wire  m_154_io_s; // @[MUL.scala 102:19]
  wire  m_154_io_cout; // @[MUL.scala 102:19]
  wire  m_155_io_x1; // @[MUL.scala 102:19]
  wire  m_155_io_x2; // @[MUL.scala 102:19]
  wire  m_155_io_x3; // @[MUL.scala 102:19]
  wire  m_155_io_s; // @[MUL.scala 102:19]
  wire  m_155_io_cout; // @[MUL.scala 102:19]
  wire  m_156_io_x1; // @[MUL.scala 102:19]
  wire  m_156_io_x2; // @[MUL.scala 102:19]
  wire  m_156_io_x3; // @[MUL.scala 102:19]
  wire  m_156_io_s; // @[MUL.scala 102:19]
  wire  m_156_io_cout; // @[MUL.scala 102:19]
  wire  m_157_io_x1; // @[MUL.scala 102:19]
  wire  m_157_io_x2; // @[MUL.scala 102:19]
  wire  m_157_io_x3; // @[MUL.scala 102:19]
  wire  m_157_io_s; // @[MUL.scala 102:19]
  wire  m_157_io_cout; // @[MUL.scala 102:19]
  wire  m_158_io_x1; // @[MUL.scala 102:19]
  wire  m_158_io_x2; // @[MUL.scala 102:19]
  wire  m_158_io_x3; // @[MUL.scala 102:19]
  wire  m_158_io_s; // @[MUL.scala 102:19]
  wire  m_158_io_cout; // @[MUL.scala 102:19]
  wire  m_159_io_x1; // @[MUL.scala 102:19]
  wire  m_159_io_x2; // @[MUL.scala 102:19]
  wire  m_159_io_x3; // @[MUL.scala 102:19]
  wire  m_159_io_s; // @[MUL.scala 102:19]
  wire  m_159_io_cout; // @[MUL.scala 102:19]
  wire  m_160_io_x1; // @[MUL.scala 102:19]
  wire  m_160_io_x2; // @[MUL.scala 102:19]
  wire  m_160_io_x3; // @[MUL.scala 102:19]
  wire  m_160_io_s; // @[MUL.scala 102:19]
  wire  m_160_io_cout; // @[MUL.scala 102:19]
  wire  m_161_io_x1; // @[MUL.scala 102:19]
  wire  m_161_io_x2; // @[MUL.scala 102:19]
  wire  m_161_io_x3; // @[MUL.scala 102:19]
  wire  m_161_io_s; // @[MUL.scala 102:19]
  wire  m_161_io_cout; // @[MUL.scala 102:19]
  wire  m_162_io_x1; // @[MUL.scala 102:19]
  wire  m_162_io_x2; // @[MUL.scala 102:19]
  wire  m_162_io_x3; // @[MUL.scala 102:19]
  wire  m_162_io_s; // @[MUL.scala 102:19]
  wire  m_162_io_cout; // @[MUL.scala 102:19]
  wire  m_163_io_x1; // @[MUL.scala 102:19]
  wire  m_163_io_x2; // @[MUL.scala 102:19]
  wire  m_163_io_x3; // @[MUL.scala 102:19]
  wire  m_163_io_s; // @[MUL.scala 102:19]
  wire  m_163_io_cout; // @[MUL.scala 102:19]
  wire  m_164_io_x1; // @[MUL.scala 102:19]
  wire  m_164_io_x2; // @[MUL.scala 102:19]
  wire  m_164_io_x3; // @[MUL.scala 102:19]
  wire  m_164_io_s; // @[MUL.scala 102:19]
  wire  m_164_io_cout; // @[MUL.scala 102:19]
  wire  m_165_io_in_0; // @[MUL.scala 124:19]
  wire  m_165_io_in_1; // @[MUL.scala 124:19]
  wire  m_165_io_out_0; // @[MUL.scala 124:19]
  wire  m_165_io_out_1; // @[MUL.scala 124:19]
  wire  m_166_io_x1; // @[MUL.scala 102:19]
  wire  m_166_io_x2; // @[MUL.scala 102:19]
  wire  m_166_io_x3; // @[MUL.scala 102:19]
  wire  m_166_io_s; // @[MUL.scala 102:19]
  wire  m_166_io_cout; // @[MUL.scala 102:19]
  wire  m_167_io_x1; // @[MUL.scala 102:19]
  wire  m_167_io_x2; // @[MUL.scala 102:19]
  wire  m_167_io_x3; // @[MUL.scala 102:19]
  wire  m_167_io_s; // @[MUL.scala 102:19]
  wire  m_167_io_cout; // @[MUL.scala 102:19]
  wire  m_168_io_x1; // @[MUL.scala 102:19]
  wire  m_168_io_x2; // @[MUL.scala 102:19]
  wire  m_168_io_x3; // @[MUL.scala 102:19]
  wire  m_168_io_s; // @[MUL.scala 102:19]
  wire  m_168_io_cout; // @[MUL.scala 102:19]
  wire  m_169_io_x1; // @[MUL.scala 102:19]
  wire  m_169_io_x2; // @[MUL.scala 102:19]
  wire  m_169_io_x3; // @[MUL.scala 102:19]
  wire  m_169_io_s; // @[MUL.scala 102:19]
  wire  m_169_io_cout; // @[MUL.scala 102:19]
  wire  m_170_io_x1; // @[MUL.scala 102:19]
  wire  m_170_io_x2; // @[MUL.scala 102:19]
  wire  m_170_io_x3; // @[MUL.scala 102:19]
  wire  m_170_io_s; // @[MUL.scala 102:19]
  wire  m_170_io_cout; // @[MUL.scala 102:19]
  wire  m_171_io_x1; // @[MUL.scala 102:19]
  wire  m_171_io_x2; // @[MUL.scala 102:19]
  wire  m_171_io_x3; // @[MUL.scala 102:19]
  wire  m_171_io_s; // @[MUL.scala 102:19]
  wire  m_171_io_cout; // @[MUL.scala 102:19]
  wire  m_172_io_in_0; // @[MUL.scala 124:19]
  wire  m_172_io_in_1; // @[MUL.scala 124:19]
  wire  m_172_io_out_0; // @[MUL.scala 124:19]
  wire  m_172_io_out_1; // @[MUL.scala 124:19]
  wire  m_173_io_x1; // @[MUL.scala 102:19]
  wire  m_173_io_x2; // @[MUL.scala 102:19]
  wire  m_173_io_x3; // @[MUL.scala 102:19]
  wire  m_173_io_s; // @[MUL.scala 102:19]
  wire  m_173_io_cout; // @[MUL.scala 102:19]
  wire  m_174_io_x1; // @[MUL.scala 102:19]
  wire  m_174_io_x2; // @[MUL.scala 102:19]
  wire  m_174_io_x3; // @[MUL.scala 102:19]
  wire  m_174_io_s; // @[MUL.scala 102:19]
  wire  m_174_io_cout; // @[MUL.scala 102:19]
  wire  m_175_io_x1; // @[MUL.scala 102:19]
  wire  m_175_io_x2; // @[MUL.scala 102:19]
  wire  m_175_io_x3; // @[MUL.scala 102:19]
  wire  m_175_io_s; // @[MUL.scala 102:19]
  wire  m_175_io_cout; // @[MUL.scala 102:19]
  wire  m_176_io_x1; // @[MUL.scala 102:19]
  wire  m_176_io_x2; // @[MUL.scala 102:19]
  wire  m_176_io_x3; // @[MUL.scala 102:19]
  wire  m_176_io_s; // @[MUL.scala 102:19]
  wire  m_176_io_cout; // @[MUL.scala 102:19]
  wire  m_177_io_x1; // @[MUL.scala 102:19]
  wire  m_177_io_x2; // @[MUL.scala 102:19]
  wire  m_177_io_x3; // @[MUL.scala 102:19]
  wire  m_177_io_s; // @[MUL.scala 102:19]
  wire  m_177_io_cout; // @[MUL.scala 102:19]
  wire  m_178_io_x1; // @[MUL.scala 102:19]
  wire  m_178_io_x2; // @[MUL.scala 102:19]
  wire  m_178_io_x3; // @[MUL.scala 102:19]
  wire  m_178_io_s; // @[MUL.scala 102:19]
  wire  m_178_io_cout; // @[MUL.scala 102:19]
  wire  m_179_io_x1; // @[MUL.scala 102:19]
  wire  m_179_io_x2; // @[MUL.scala 102:19]
  wire  m_179_io_x3; // @[MUL.scala 102:19]
  wire  m_179_io_s; // @[MUL.scala 102:19]
  wire  m_179_io_cout; // @[MUL.scala 102:19]
  wire  m_180_io_x1; // @[MUL.scala 102:19]
  wire  m_180_io_x2; // @[MUL.scala 102:19]
  wire  m_180_io_x3; // @[MUL.scala 102:19]
  wire  m_180_io_s; // @[MUL.scala 102:19]
  wire  m_180_io_cout; // @[MUL.scala 102:19]
  wire  m_181_io_x1; // @[MUL.scala 102:19]
  wire  m_181_io_x2; // @[MUL.scala 102:19]
  wire  m_181_io_x3; // @[MUL.scala 102:19]
  wire  m_181_io_s; // @[MUL.scala 102:19]
  wire  m_181_io_cout; // @[MUL.scala 102:19]
  wire  m_182_io_x1; // @[MUL.scala 102:19]
  wire  m_182_io_x2; // @[MUL.scala 102:19]
  wire  m_182_io_x3; // @[MUL.scala 102:19]
  wire  m_182_io_s; // @[MUL.scala 102:19]
  wire  m_182_io_cout; // @[MUL.scala 102:19]
  wire  m_183_io_x1; // @[MUL.scala 102:19]
  wire  m_183_io_x2; // @[MUL.scala 102:19]
  wire  m_183_io_x3; // @[MUL.scala 102:19]
  wire  m_183_io_s; // @[MUL.scala 102:19]
  wire  m_183_io_cout; // @[MUL.scala 102:19]
  wire  m_184_io_x1; // @[MUL.scala 102:19]
  wire  m_184_io_x2; // @[MUL.scala 102:19]
  wire  m_184_io_x3; // @[MUL.scala 102:19]
  wire  m_184_io_s; // @[MUL.scala 102:19]
  wire  m_184_io_cout; // @[MUL.scala 102:19]
  wire  m_185_io_x1; // @[MUL.scala 102:19]
  wire  m_185_io_x2; // @[MUL.scala 102:19]
  wire  m_185_io_x3; // @[MUL.scala 102:19]
  wire  m_185_io_s; // @[MUL.scala 102:19]
  wire  m_185_io_cout; // @[MUL.scala 102:19]
  wire  m_186_io_x1; // @[MUL.scala 102:19]
  wire  m_186_io_x2; // @[MUL.scala 102:19]
  wire  m_186_io_x3; // @[MUL.scala 102:19]
  wire  m_186_io_s; // @[MUL.scala 102:19]
  wire  m_186_io_cout; // @[MUL.scala 102:19]
  wire  m_187_io_x1; // @[MUL.scala 102:19]
  wire  m_187_io_x2; // @[MUL.scala 102:19]
  wire  m_187_io_x3; // @[MUL.scala 102:19]
  wire  m_187_io_s; // @[MUL.scala 102:19]
  wire  m_187_io_cout; // @[MUL.scala 102:19]
  wire  m_188_io_x1; // @[MUL.scala 102:19]
  wire  m_188_io_x2; // @[MUL.scala 102:19]
  wire  m_188_io_x3; // @[MUL.scala 102:19]
  wire  m_188_io_s; // @[MUL.scala 102:19]
  wire  m_188_io_cout; // @[MUL.scala 102:19]
  wire  m_189_io_x1; // @[MUL.scala 102:19]
  wire  m_189_io_x2; // @[MUL.scala 102:19]
  wire  m_189_io_x3; // @[MUL.scala 102:19]
  wire  m_189_io_s; // @[MUL.scala 102:19]
  wire  m_189_io_cout; // @[MUL.scala 102:19]
  wire  m_190_io_x1; // @[MUL.scala 102:19]
  wire  m_190_io_x2; // @[MUL.scala 102:19]
  wire  m_190_io_x3; // @[MUL.scala 102:19]
  wire  m_190_io_s; // @[MUL.scala 102:19]
  wire  m_190_io_cout; // @[MUL.scala 102:19]
  wire  m_191_io_x1; // @[MUL.scala 102:19]
  wire  m_191_io_x2; // @[MUL.scala 102:19]
  wire  m_191_io_x3; // @[MUL.scala 102:19]
  wire  m_191_io_s; // @[MUL.scala 102:19]
  wire  m_191_io_cout; // @[MUL.scala 102:19]
  wire  m_192_io_x1; // @[MUL.scala 102:19]
  wire  m_192_io_x2; // @[MUL.scala 102:19]
  wire  m_192_io_x3; // @[MUL.scala 102:19]
  wire  m_192_io_s; // @[MUL.scala 102:19]
  wire  m_192_io_cout; // @[MUL.scala 102:19]
  wire  m_193_io_x1; // @[MUL.scala 102:19]
  wire  m_193_io_x2; // @[MUL.scala 102:19]
  wire  m_193_io_x3; // @[MUL.scala 102:19]
  wire  m_193_io_s; // @[MUL.scala 102:19]
  wire  m_193_io_cout; // @[MUL.scala 102:19]
  wire  m_194_io_x1; // @[MUL.scala 102:19]
  wire  m_194_io_x2; // @[MUL.scala 102:19]
  wire  m_194_io_x3; // @[MUL.scala 102:19]
  wire  m_194_io_s; // @[MUL.scala 102:19]
  wire  m_194_io_cout; // @[MUL.scala 102:19]
  wire  m_195_io_x1; // @[MUL.scala 102:19]
  wire  m_195_io_x2; // @[MUL.scala 102:19]
  wire  m_195_io_x3; // @[MUL.scala 102:19]
  wire  m_195_io_s; // @[MUL.scala 102:19]
  wire  m_195_io_cout; // @[MUL.scala 102:19]
  wire  m_196_io_x1; // @[MUL.scala 102:19]
  wire  m_196_io_x2; // @[MUL.scala 102:19]
  wire  m_196_io_x3; // @[MUL.scala 102:19]
  wire  m_196_io_s; // @[MUL.scala 102:19]
  wire  m_196_io_cout; // @[MUL.scala 102:19]
  wire  m_197_io_x1; // @[MUL.scala 102:19]
  wire  m_197_io_x2; // @[MUL.scala 102:19]
  wire  m_197_io_x3; // @[MUL.scala 102:19]
  wire  m_197_io_s; // @[MUL.scala 102:19]
  wire  m_197_io_cout; // @[MUL.scala 102:19]
  wire  m_198_io_x1; // @[MUL.scala 102:19]
  wire  m_198_io_x2; // @[MUL.scala 102:19]
  wire  m_198_io_x3; // @[MUL.scala 102:19]
  wire  m_198_io_s; // @[MUL.scala 102:19]
  wire  m_198_io_cout; // @[MUL.scala 102:19]
  wire  m_199_io_x1; // @[MUL.scala 102:19]
  wire  m_199_io_x2; // @[MUL.scala 102:19]
  wire  m_199_io_x3; // @[MUL.scala 102:19]
  wire  m_199_io_s; // @[MUL.scala 102:19]
  wire  m_199_io_cout; // @[MUL.scala 102:19]
  wire  m_200_io_x1; // @[MUL.scala 102:19]
  wire  m_200_io_x2; // @[MUL.scala 102:19]
  wire  m_200_io_x3; // @[MUL.scala 102:19]
  wire  m_200_io_s; // @[MUL.scala 102:19]
  wire  m_200_io_cout; // @[MUL.scala 102:19]
  wire  m_201_io_x1; // @[MUL.scala 102:19]
  wire  m_201_io_x2; // @[MUL.scala 102:19]
  wire  m_201_io_x3; // @[MUL.scala 102:19]
  wire  m_201_io_s; // @[MUL.scala 102:19]
  wire  m_201_io_cout; // @[MUL.scala 102:19]
  wire  m_202_io_x1; // @[MUL.scala 102:19]
  wire  m_202_io_x2; // @[MUL.scala 102:19]
  wire  m_202_io_x3; // @[MUL.scala 102:19]
  wire  m_202_io_s; // @[MUL.scala 102:19]
  wire  m_202_io_cout; // @[MUL.scala 102:19]
  wire  m_203_io_x1; // @[MUL.scala 102:19]
  wire  m_203_io_x2; // @[MUL.scala 102:19]
  wire  m_203_io_x3; // @[MUL.scala 102:19]
  wire  m_203_io_s; // @[MUL.scala 102:19]
  wire  m_203_io_cout; // @[MUL.scala 102:19]
  wire  m_204_io_x1; // @[MUL.scala 102:19]
  wire  m_204_io_x2; // @[MUL.scala 102:19]
  wire  m_204_io_x3; // @[MUL.scala 102:19]
  wire  m_204_io_s; // @[MUL.scala 102:19]
  wire  m_204_io_cout; // @[MUL.scala 102:19]
  wire  m_205_io_x1; // @[MUL.scala 102:19]
  wire  m_205_io_x2; // @[MUL.scala 102:19]
  wire  m_205_io_x3; // @[MUL.scala 102:19]
  wire  m_205_io_s; // @[MUL.scala 102:19]
  wire  m_205_io_cout; // @[MUL.scala 102:19]
  wire  m_206_io_x1; // @[MUL.scala 102:19]
  wire  m_206_io_x2; // @[MUL.scala 102:19]
  wire  m_206_io_x3; // @[MUL.scala 102:19]
  wire  m_206_io_s; // @[MUL.scala 102:19]
  wire  m_206_io_cout; // @[MUL.scala 102:19]
  wire  m_207_io_x1; // @[MUL.scala 102:19]
  wire  m_207_io_x2; // @[MUL.scala 102:19]
  wire  m_207_io_x3; // @[MUL.scala 102:19]
  wire  m_207_io_s; // @[MUL.scala 102:19]
  wire  m_207_io_cout; // @[MUL.scala 102:19]
  wire  m_208_io_in_0; // @[MUL.scala 124:19]
  wire  m_208_io_in_1; // @[MUL.scala 124:19]
  wire  m_208_io_out_0; // @[MUL.scala 124:19]
  wire  m_208_io_out_1; // @[MUL.scala 124:19]
  wire  m_209_io_x1; // @[MUL.scala 102:19]
  wire  m_209_io_x2; // @[MUL.scala 102:19]
  wire  m_209_io_x3; // @[MUL.scala 102:19]
  wire  m_209_io_s; // @[MUL.scala 102:19]
  wire  m_209_io_cout; // @[MUL.scala 102:19]
  wire  m_210_io_x1; // @[MUL.scala 102:19]
  wire  m_210_io_x2; // @[MUL.scala 102:19]
  wire  m_210_io_x3; // @[MUL.scala 102:19]
  wire  m_210_io_s; // @[MUL.scala 102:19]
  wire  m_210_io_cout; // @[MUL.scala 102:19]
  wire  m_211_io_x1; // @[MUL.scala 102:19]
  wire  m_211_io_x2; // @[MUL.scala 102:19]
  wire  m_211_io_x3; // @[MUL.scala 102:19]
  wire  m_211_io_s; // @[MUL.scala 102:19]
  wire  m_211_io_cout; // @[MUL.scala 102:19]
  wire  m_212_io_x1; // @[MUL.scala 102:19]
  wire  m_212_io_x2; // @[MUL.scala 102:19]
  wire  m_212_io_x3; // @[MUL.scala 102:19]
  wire  m_212_io_s; // @[MUL.scala 102:19]
  wire  m_212_io_cout; // @[MUL.scala 102:19]
  wire  m_213_io_x1; // @[MUL.scala 102:19]
  wire  m_213_io_x2; // @[MUL.scala 102:19]
  wire  m_213_io_x3; // @[MUL.scala 102:19]
  wire  m_213_io_s; // @[MUL.scala 102:19]
  wire  m_213_io_cout; // @[MUL.scala 102:19]
  wire  m_214_io_x1; // @[MUL.scala 102:19]
  wire  m_214_io_x2; // @[MUL.scala 102:19]
  wire  m_214_io_x3; // @[MUL.scala 102:19]
  wire  m_214_io_s; // @[MUL.scala 102:19]
  wire  m_214_io_cout; // @[MUL.scala 102:19]
  wire  m_215_io_x1; // @[MUL.scala 102:19]
  wire  m_215_io_x2; // @[MUL.scala 102:19]
  wire  m_215_io_x3; // @[MUL.scala 102:19]
  wire  m_215_io_s; // @[MUL.scala 102:19]
  wire  m_215_io_cout; // @[MUL.scala 102:19]
  wire  m_216_io_in_0; // @[MUL.scala 124:19]
  wire  m_216_io_in_1; // @[MUL.scala 124:19]
  wire  m_216_io_out_0; // @[MUL.scala 124:19]
  wire  m_216_io_out_1; // @[MUL.scala 124:19]
  wire  m_217_io_x1; // @[MUL.scala 102:19]
  wire  m_217_io_x2; // @[MUL.scala 102:19]
  wire  m_217_io_x3; // @[MUL.scala 102:19]
  wire  m_217_io_s; // @[MUL.scala 102:19]
  wire  m_217_io_cout; // @[MUL.scala 102:19]
  wire  m_218_io_x1; // @[MUL.scala 102:19]
  wire  m_218_io_x2; // @[MUL.scala 102:19]
  wire  m_218_io_x3; // @[MUL.scala 102:19]
  wire  m_218_io_s; // @[MUL.scala 102:19]
  wire  m_218_io_cout; // @[MUL.scala 102:19]
  wire  m_219_io_x1; // @[MUL.scala 102:19]
  wire  m_219_io_x2; // @[MUL.scala 102:19]
  wire  m_219_io_x3; // @[MUL.scala 102:19]
  wire  m_219_io_s; // @[MUL.scala 102:19]
  wire  m_219_io_cout; // @[MUL.scala 102:19]
  wire  m_220_io_x1; // @[MUL.scala 102:19]
  wire  m_220_io_x2; // @[MUL.scala 102:19]
  wire  m_220_io_x3; // @[MUL.scala 102:19]
  wire  m_220_io_s; // @[MUL.scala 102:19]
  wire  m_220_io_cout; // @[MUL.scala 102:19]
  wire  m_221_io_x1; // @[MUL.scala 102:19]
  wire  m_221_io_x2; // @[MUL.scala 102:19]
  wire  m_221_io_x3; // @[MUL.scala 102:19]
  wire  m_221_io_s; // @[MUL.scala 102:19]
  wire  m_221_io_cout; // @[MUL.scala 102:19]
  wire  m_222_io_x1; // @[MUL.scala 102:19]
  wire  m_222_io_x2; // @[MUL.scala 102:19]
  wire  m_222_io_x3; // @[MUL.scala 102:19]
  wire  m_222_io_s; // @[MUL.scala 102:19]
  wire  m_222_io_cout; // @[MUL.scala 102:19]
  wire  m_223_io_x1; // @[MUL.scala 102:19]
  wire  m_223_io_x2; // @[MUL.scala 102:19]
  wire  m_223_io_x3; // @[MUL.scala 102:19]
  wire  m_223_io_s; // @[MUL.scala 102:19]
  wire  m_223_io_cout; // @[MUL.scala 102:19]
  wire  m_224_io_x1; // @[MUL.scala 102:19]
  wire  m_224_io_x2; // @[MUL.scala 102:19]
  wire  m_224_io_x3; // @[MUL.scala 102:19]
  wire  m_224_io_s; // @[MUL.scala 102:19]
  wire  m_224_io_cout; // @[MUL.scala 102:19]
  wire  m_225_io_x1; // @[MUL.scala 102:19]
  wire  m_225_io_x2; // @[MUL.scala 102:19]
  wire  m_225_io_x3; // @[MUL.scala 102:19]
  wire  m_225_io_s; // @[MUL.scala 102:19]
  wire  m_225_io_cout; // @[MUL.scala 102:19]
  wire  m_226_io_x1; // @[MUL.scala 102:19]
  wire  m_226_io_x2; // @[MUL.scala 102:19]
  wire  m_226_io_x3; // @[MUL.scala 102:19]
  wire  m_226_io_s; // @[MUL.scala 102:19]
  wire  m_226_io_cout; // @[MUL.scala 102:19]
  wire  m_227_io_x1; // @[MUL.scala 102:19]
  wire  m_227_io_x2; // @[MUL.scala 102:19]
  wire  m_227_io_x3; // @[MUL.scala 102:19]
  wire  m_227_io_s; // @[MUL.scala 102:19]
  wire  m_227_io_cout; // @[MUL.scala 102:19]
  wire  m_228_io_x1; // @[MUL.scala 102:19]
  wire  m_228_io_x2; // @[MUL.scala 102:19]
  wire  m_228_io_x3; // @[MUL.scala 102:19]
  wire  m_228_io_s; // @[MUL.scala 102:19]
  wire  m_228_io_cout; // @[MUL.scala 102:19]
  wire  m_229_io_x1; // @[MUL.scala 102:19]
  wire  m_229_io_x2; // @[MUL.scala 102:19]
  wire  m_229_io_x3; // @[MUL.scala 102:19]
  wire  m_229_io_s; // @[MUL.scala 102:19]
  wire  m_229_io_cout; // @[MUL.scala 102:19]
  wire  m_230_io_x1; // @[MUL.scala 102:19]
  wire  m_230_io_x2; // @[MUL.scala 102:19]
  wire  m_230_io_x3; // @[MUL.scala 102:19]
  wire  m_230_io_s; // @[MUL.scala 102:19]
  wire  m_230_io_cout; // @[MUL.scala 102:19]
  wire  m_231_io_x1; // @[MUL.scala 102:19]
  wire  m_231_io_x2; // @[MUL.scala 102:19]
  wire  m_231_io_x3; // @[MUL.scala 102:19]
  wire  m_231_io_s; // @[MUL.scala 102:19]
  wire  m_231_io_cout; // @[MUL.scala 102:19]
  wire  m_232_io_x1; // @[MUL.scala 102:19]
  wire  m_232_io_x2; // @[MUL.scala 102:19]
  wire  m_232_io_x3; // @[MUL.scala 102:19]
  wire  m_232_io_s; // @[MUL.scala 102:19]
  wire  m_232_io_cout; // @[MUL.scala 102:19]
  wire  m_233_io_x1; // @[MUL.scala 102:19]
  wire  m_233_io_x2; // @[MUL.scala 102:19]
  wire  m_233_io_x3; // @[MUL.scala 102:19]
  wire  m_233_io_s; // @[MUL.scala 102:19]
  wire  m_233_io_cout; // @[MUL.scala 102:19]
  wire  m_234_io_x1; // @[MUL.scala 102:19]
  wire  m_234_io_x2; // @[MUL.scala 102:19]
  wire  m_234_io_x3; // @[MUL.scala 102:19]
  wire  m_234_io_s; // @[MUL.scala 102:19]
  wire  m_234_io_cout; // @[MUL.scala 102:19]
  wire  m_235_io_x1; // @[MUL.scala 102:19]
  wire  m_235_io_x2; // @[MUL.scala 102:19]
  wire  m_235_io_x3; // @[MUL.scala 102:19]
  wire  m_235_io_s; // @[MUL.scala 102:19]
  wire  m_235_io_cout; // @[MUL.scala 102:19]
  wire  m_236_io_x1; // @[MUL.scala 102:19]
  wire  m_236_io_x2; // @[MUL.scala 102:19]
  wire  m_236_io_x3; // @[MUL.scala 102:19]
  wire  m_236_io_s; // @[MUL.scala 102:19]
  wire  m_236_io_cout; // @[MUL.scala 102:19]
  wire  m_237_io_x1; // @[MUL.scala 102:19]
  wire  m_237_io_x2; // @[MUL.scala 102:19]
  wire  m_237_io_x3; // @[MUL.scala 102:19]
  wire  m_237_io_s; // @[MUL.scala 102:19]
  wire  m_237_io_cout; // @[MUL.scala 102:19]
  wire  m_238_io_x1; // @[MUL.scala 102:19]
  wire  m_238_io_x2; // @[MUL.scala 102:19]
  wire  m_238_io_x3; // @[MUL.scala 102:19]
  wire  m_238_io_s; // @[MUL.scala 102:19]
  wire  m_238_io_cout; // @[MUL.scala 102:19]
  wire  m_239_io_x1; // @[MUL.scala 102:19]
  wire  m_239_io_x2; // @[MUL.scala 102:19]
  wire  m_239_io_x3; // @[MUL.scala 102:19]
  wire  m_239_io_s; // @[MUL.scala 102:19]
  wire  m_239_io_cout; // @[MUL.scala 102:19]
  wire  m_240_io_x1; // @[MUL.scala 102:19]
  wire  m_240_io_x2; // @[MUL.scala 102:19]
  wire  m_240_io_x3; // @[MUL.scala 102:19]
  wire  m_240_io_s; // @[MUL.scala 102:19]
  wire  m_240_io_cout; // @[MUL.scala 102:19]
  wire  m_241_io_x1; // @[MUL.scala 102:19]
  wire  m_241_io_x2; // @[MUL.scala 102:19]
  wire  m_241_io_x3; // @[MUL.scala 102:19]
  wire  m_241_io_s; // @[MUL.scala 102:19]
  wire  m_241_io_cout; // @[MUL.scala 102:19]
  wire  m_242_io_x1; // @[MUL.scala 102:19]
  wire  m_242_io_x2; // @[MUL.scala 102:19]
  wire  m_242_io_x3; // @[MUL.scala 102:19]
  wire  m_242_io_s; // @[MUL.scala 102:19]
  wire  m_242_io_cout; // @[MUL.scala 102:19]
  wire  m_243_io_x1; // @[MUL.scala 102:19]
  wire  m_243_io_x2; // @[MUL.scala 102:19]
  wire  m_243_io_x3; // @[MUL.scala 102:19]
  wire  m_243_io_s; // @[MUL.scala 102:19]
  wire  m_243_io_cout; // @[MUL.scala 102:19]
  wire  m_244_io_x1; // @[MUL.scala 102:19]
  wire  m_244_io_x2; // @[MUL.scala 102:19]
  wire  m_244_io_x3; // @[MUL.scala 102:19]
  wire  m_244_io_s; // @[MUL.scala 102:19]
  wire  m_244_io_cout; // @[MUL.scala 102:19]
  wire  m_245_io_x1; // @[MUL.scala 102:19]
  wire  m_245_io_x2; // @[MUL.scala 102:19]
  wire  m_245_io_x3; // @[MUL.scala 102:19]
  wire  m_245_io_s; // @[MUL.scala 102:19]
  wire  m_245_io_cout; // @[MUL.scala 102:19]
  wire  m_246_io_x1; // @[MUL.scala 102:19]
  wire  m_246_io_x2; // @[MUL.scala 102:19]
  wire  m_246_io_x3; // @[MUL.scala 102:19]
  wire  m_246_io_s; // @[MUL.scala 102:19]
  wire  m_246_io_cout; // @[MUL.scala 102:19]
  wire  m_247_io_x1; // @[MUL.scala 102:19]
  wire  m_247_io_x2; // @[MUL.scala 102:19]
  wire  m_247_io_x3; // @[MUL.scala 102:19]
  wire  m_247_io_s; // @[MUL.scala 102:19]
  wire  m_247_io_cout; // @[MUL.scala 102:19]
  wire  m_248_io_x1; // @[MUL.scala 102:19]
  wire  m_248_io_x2; // @[MUL.scala 102:19]
  wire  m_248_io_x3; // @[MUL.scala 102:19]
  wire  m_248_io_s; // @[MUL.scala 102:19]
  wire  m_248_io_cout; // @[MUL.scala 102:19]
  wire  m_249_io_x1; // @[MUL.scala 102:19]
  wire  m_249_io_x2; // @[MUL.scala 102:19]
  wire  m_249_io_x3; // @[MUL.scala 102:19]
  wire  m_249_io_s; // @[MUL.scala 102:19]
  wire  m_249_io_cout; // @[MUL.scala 102:19]
  wire  m_250_io_x1; // @[MUL.scala 102:19]
  wire  m_250_io_x2; // @[MUL.scala 102:19]
  wire  m_250_io_x3; // @[MUL.scala 102:19]
  wire  m_250_io_s; // @[MUL.scala 102:19]
  wire  m_250_io_cout; // @[MUL.scala 102:19]
  wire  m_251_io_x1; // @[MUL.scala 102:19]
  wire  m_251_io_x2; // @[MUL.scala 102:19]
  wire  m_251_io_x3; // @[MUL.scala 102:19]
  wire  m_251_io_s; // @[MUL.scala 102:19]
  wire  m_251_io_cout; // @[MUL.scala 102:19]
  wire  m_252_io_x1; // @[MUL.scala 102:19]
  wire  m_252_io_x2; // @[MUL.scala 102:19]
  wire  m_252_io_x3; // @[MUL.scala 102:19]
  wire  m_252_io_s; // @[MUL.scala 102:19]
  wire  m_252_io_cout; // @[MUL.scala 102:19]
  wire  m_253_io_x1; // @[MUL.scala 102:19]
  wire  m_253_io_x2; // @[MUL.scala 102:19]
  wire  m_253_io_x3; // @[MUL.scala 102:19]
  wire  m_253_io_s; // @[MUL.scala 102:19]
  wire  m_253_io_cout; // @[MUL.scala 102:19]
  wire  m_254_io_x1; // @[MUL.scala 102:19]
  wire  m_254_io_x2; // @[MUL.scala 102:19]
  wire  m_254_io_x3; // @[MUL.scala 102:19]
  wire  m_254_io_s; // @[MUL.scala 102:19]
  wire  m_254_io_cout; // @[MUL.scala 102:19]
  wire  m_255_io_x1; // @[MUL.scala 102:19]
  wire  m_255_io_x2; // @[MUL.scala 102:19]
  wire  m_255_io_x3; // @[MUL.scala 102:19]
  wire  m_255_io_s; // @[MUL.scala 102:19]
  wire  m_255_io_cout; // @[MUL.scala 102:19]
  wire  m_256_io_x1; // @[MUL.scala 102:19]
  wire  m_256_io_x2; // @[MUL.scala 102:19]
  wire  m_256_io_x3; // @[MUL.scala 102:19]
  wire  m_256_io_s; // @[MUL.scala 102:19]
  wire  m_256_io_cout; // @[MUL.scala 102:19]
  wire  m_257_io_in_0; // @[MUL.scala 124:19]
  wire  m_257_io_in_1; // @[MUL.scala 124:19]
  wire  m_257_io_out_0; // @[MUL.scala 124:19]
  wire  m_257_io_out_1; // @[MUL.scala 124:19]
  wire  m_258_io_x1; // @[MUL.scala 102:19]
  wire  m_258_io_x2; // @[MUL.scala 102:19]
  wire  m_258_io_x3; // @[MUL.scala 102:19]
  wire  m_258_io_s; // @[MUL.scala 102:19]
  wire  m_258_io_cout; // @[MUL.scala 102:19]
  wire  m_259_io_x1; // @[MUL.scala 102:19]
  wire  m_259_io_x2; // @[MUL.scala 102:19]
  wire  m_259_io_x3; // @[MUL.scala 102:19]
  wire  m_259_io_s; // @[MUL.scala 102:19]
  wire  m_259_io_cout; // @[MUL.scala 102:19]
  wire  m_260_io_x1; // @[MUL.scala 102:19]
  wire  m_260_io_x2; // @[MUL.scala 102:19]
  wire  m_260_io_x3; // @[MUL.scala 102:19]
  wire  m_260_io_s; // @[MUL.scala 102:19]
  wire  m_260_io_cout; // @[MUL.scala 102:19]
  wire  m_261_io_x1; // @[MUL.scala 102:19]
  wire  m_261_io_x2; // @[MUL.scala 102:19]
  wire  m_261_io_x3; // @[MUL.scala 102:19]
  wire  m_261_io_s; // @[MUL.scala 102:19]
  wire  m_261_io_cout; // @[MUL.scala 102:19]
  wire  m_262_io_x1; // @[MUL.scala 102:19]
  wire  m_262_io_x2; // @[MUL.scala 102:19]
  wire  m_262_io_x3; // @[MUL.scala 102:19]
  wire  m_262_io_s; // @[MUL.scala 102:19]
  wire  m_262_io_cout; // @[MUL.scala 102:19]
  wire  m_263_io_x1; // @[MUL.scala 102:19]
  wire  m_263_io_x2; // @[MUL.scala 102:19]
  wire  m_263_io_x3; // @[MUL.scala 102:19]
  wire  m_263_io_s; // @[MUL.scala 102:19]
  wire  m_263_io_cout; // @[MUL.scala 102:19]
  wire  m_264_io_x1; // @[MUL.scala 102:19]
  wire  m_264_io_x2; // @[MUL.scala 102:19]
  wire  m_264_io_x3; // @[MUL.scala 102:19]
  wire  m_264_io_s; // @[MUL.scala 102:19]
  wire  m_264_io_cout; // @[MUL.scala 102:19]
  wire  m_265_io_x1; // @[MUL.scala 102:19]
  wire  m_265_io_x2; // @[MUL.scala 102:19]
  wire  m_265_io_x3; // @[MUL.scala 102:19]
  wire  m_265_io_s; // @[MUL.scala 102:19]
  wire  m_265_io_cout; // @[MUL.scala 102:19]
  wire  m_266_io_in_0; // @[MUL.scala 124:19]
  wire  m_266_io_in_1; // @[MUL.scala 124:19]
  wire  m_266_io_out_0; // @[MUL.scala 124:19]
  wire  m_266_io_out_1; // @[MUL.scala 124:19]
  wire  m_267_io_x1; // @[MUL.scala 102:19]
  wire  m_267_io_x2; // @[MUL.scala 102:19]
  wire  m_267_io_x3; // @[MUL.scala 102:19]
  wire  m_267_io_s; // @[MUL.scala 102:19]
  wire  m_267_io_cout; // @[MUL.scala 102:19]
  wire  m_268_io_x1; // @[MUL.scala 102:19]
  wire  m_268_io_x2; // @[MUL.scala 102:19]
  wire  m_268_io_x3; // @[MUL.scala 102:19]
  wire  m_268_io_s; // @[MUL.scala 102:19]
  wire  m_268_io_cout; // @[MUL.scala 102:19]
  wire  m_269_io_x1; // @[MUL.scala 102:19]
  wire  m_269_io_x2; // @[MUL.scala 102:19]
  wire  m_269_io_x3; // @[MUL.scala 102:19]
  wire  m_269_io_s; // @[MUL.scala 102:19]
  wire  m_269_io_cout; // @[MUL.scala 102:19]
  wire  m_270_io_x1; // @[MUL.scala 102:19]
  wire  m_270_io_x2; // @[MUL.scala 102:19]
  wire  m_270_io_x3; // @[MUL.scala 102:19]
  wire  m_270_io_s; // @[MUL.scala 102:19]
  wire  m_270_io_cout; // @[MUL.scala 102:19]
  wire  m_271_io_x1; // @[MUL.scala 102:19]
  wire  m_271_io_x2; // @[MUL.scala 102:19]
  wire  m_271_io_x3; // @[MUL.scala 102:19]
  wire  m_271_io_s; // @[MUL.scala 102:19]
  wire  m_271_io_cout; // @[MUL.scala 102:19]
  wire  m_272_io_x1; // @[MUL.scala 102:19]
  wire  m_272_io_x2; // @[MUL.scala 102:19]
  wire  m_272_io_x3; // @[MUL.scala 102:19]
  wire  m_272_io_s; // @[MUL.scala 102:19]
  wire  m_272_io_cout; // @[MUL.scala 102:19]
  wire  m_273_io_x1; // @[MUL.scala 102:19]
  wire  m_273_io_x2; // @[MUL.scala 102:19]
  wire  m_273_io_x3; // @[MUL.scala 102:19]
  wire  m_273_io_s; // @[MUL.scala 102:19]
  wire  m_273_io_cout; // @[MUL.scala 102:19]
  wire  m_274_io_x1; // @[MUL.scala 102:19]
  wire  m_274_io_x2; // @[MUL.scala 102:19]
  wire  m_274_io_x3; // @[MUL.scala 102:19]
  wire  m_274_io_s; // @[MUL.scala 102:19]
  wire  m_274_io_cout; // @[MUL.scala 102:19]
  wire  m_275_io_x1; // @[MUL.scala 102:19]
  wire  m_275_io_x2; // @[MUL.scala 102:19]
  wire  m_275_io_x3; // @[MUL.scala 102:19]
  wire  m_275_io_s; // @[MUL.scala 102:19]
  wire  m_275_io_cout; // @[MUL.scala 102:19]
  wire  m_276_io_x1; // @[MUL.scala 102:19]
  wire  m_276_io_x2; // @[MUL.scala 102:19]
  wire  m_276_io_x3; // @[MUL.scala 102:19]
  wire  m_276_io_s; // @[MUL.scala 102:19]
  wire  m_276_io_cout; // @[MUL.scala 102:19]
  wire  m_277_io_x1; // @[MUL.scala 102:19]
  wire  m_277_io_x2; // @[MUL.scala 102:19]
  wire  m_277_io_x3; // @[MUL.scala 102:19]
  wire  m_277_io_s; // @[MUL.scala 102:19]
  wire  m_277_io_cout; // @[MUL.scala 102:19]
  wire  m_278_io_x1; // @[MUL.scala 102:19]
  wire  m_278_io_x2; // @[MUL.scala 102:19]
  wire  m_278_io_x3; // @[MUL.scala 102:19]
  wire  m_278_io_s; // @[MUL.scala 102:19]
  wire  m_278_io_cout; // @[MUL.scala 102:19]
  wire  m_279_io_x1; // @[MUL.scala 102:19]
  wire  m_279_io_x2; // @[MUL.scala 102:19]
  wire  m_279_io_x3; // @[MUL.scala 102:19]
  wire  m_279_io_s; // @[MUL.scala 102:19]
  wire  m_279_io_cout; // @[MUL.scala 102:19]
  wire  m_280_io_x1; // @[MUL.scala 102:19]
  wire  m_280_io_x2; // @[MUL.scala 102:19]
  wire  m_280_io_x3; // @[MUL.scala 102:19]
  wire  m_280_io_s; // @[MUL.scala 102:19]
  wire  m_280_io_cout; // @[MUL.scala 102:19]
  wire  m_281_io_x1; // @[MUL.scala 102:19]
  wire  m_281_io_x2; // @[MUL.scala 102:19]
  wire  m_281_io_x3; // @[MUL.scala 102:19]
  wire  m_281_io_s; // @[MUL.scala 102:19]
  wire  m_281_io_cout; // @[MUL.scala 102:19]
  wire  m_282_io_x1; // @[MUL.scala 102:19]
  wire  m_282_io_x2; // @[MUL.scala 102:19]
  wire  m_282_io_x3; // @[MUL.scala 102:19]
  wire  m_282_io_s; // @[MUL.scala 102:19]
  wire  m_282_io_cout; // @[MUL.scala 102:19]
  wire  m_283_io_x1; // @[MUL.scala 102:19]
  wire  m_283_io_x2; // @[MUL.scala 102:19]
  wire  m_283_io_x3; // @[MUL.scala 102:19]
  wire  m_283_io_s; // @[MUL.scala 102:19]
  wire  m_283_io_cout; // @[MUL.scala 102:19]
  wire  m_284_io_x1; // @[MUL.scala 102:19]
  wire  m_284_io_x2; // @[MUL.scala 102:19]
  wire  m_284_io_x3; // @[MUL.scala 102:19]
  wire  m_284_io_s; // @[MUL.scala 102:19]
  wire  m_284_io_cout; // @[MUL.scala 102:19]
  wire  m_285_io_x1; // @[MUL.scala 102:19]
  wire  m_285_io_x2; // @[MUL.scala 102:19]
  wire  m_285_io_x3; // @[MUL.scala 102:19]
  wire  m_285_io_s; // @[MUL.scala 102:19]
  wire  m_285_io_cout; // @[MUL.scala 102:19]
  wire  m_286_io_x1; // @[MUL.scala 102:19]
  wire  m_286_io_x2; // @[MUL.scala 102:19]
  wire  m_286_io_x3; // @[MUL.scala 102:19]
  wire  m_286_io_s; // @[MUL.scala 102:19]
  wire  m_286_io_cout; // @[MUL.scala 102:19]
  wire  m_287_io_x1; // @[MUL.scala 102:19]
  wire  m_287_io_x2; // @[MUL.scala 102:19]
  wire  m_287_io_x3; // @[MUL.scala 102:19]
  wire  m_287_io_s; // @[MUL.scala 102:19]
  wire  m_287_io_cout; // @[MUL.scala 102:19]
  wire  m_288_io_x1; // @[MUL.scala 102:19]
  wire  m_288_io_x2; // @[MUL.scala 102:19]
  wire  m_288_io_x3; // @[MUL.scala 102:19]
  wire  m_288_io_s; // @[MUL.scala 102:19]
  wire  m_288_io_cout; // @[MUL.scala 102:19]
  wire  m_289_io_x1; // @[MUL.scala 102:19]
  wire  m_289_io_x2; // @[MUL.scala 102:19]
  wire  m_289_io_x3; // @[MUL.scala 102:19]
  wire  m_289_io_s; // @[MUL.scala 102:19]
  wire  m_289_io_cout; // @[MUL.scala 102:19]
  wire  m_290_io_x1; // @[MUL.scala 102:19]
  wire  m_290_io_x2; // @[MUL.scala 102:19]
  wire  m_290_io_x3; // @[MUL.scala 102:19]
  wire  m_290_io_s; // @[MUL.scala 102:19]
  wire  m_290_io_cout; // @[MUL.scala 102:19]
  wire  m_291_io_x1; // @[MUL.scala 102:19]
  wire  m_291_io_x2; // @[MUL.scala 102:19]
  wire  m_291_io_x3; // @[MUL.scala 102:19]
  wire  m_291_io_s; // @[MUL.scala 102:19]
  wire  m_291_io_cout; // @[MUL.scala 102:19]
  wire  m_292_io_x1; // @[MUL.scala 102:19]
  wire  m_292_io_x2; // @[MUL.scala 102:19]
  wire  m_292_io_x3; // @[MUL.scala 102:19]
  wire  m_292_io_s; // @[MUL.scala 102:19]
  wire  m_292_io_cout; // @[MUL.scala 102:19]
  wire  m_293_io_x1; // @[MUL.scala 102:19]
  wire  m_293_io_x2; // @[MUL.scala 102:19]
  wire  m_293_io_x3; // @[MUL.scala 102:19]
  wire  m_293_io_s; // @[MUL.scala 102:19]
  wire  m_293_io_cout; // @[MUL.scala 102:19]
  wire  m_294_io_x1; // @[MUL.scala 102:19]
  wire  m_294_io_x2; // @[MUL.scala 102:19]
  wire  m_294_io_x3; // @[MUL.scala 102:19]
  wire  m_294_io_s; // @[MUL.scala 102:19]
  wire  m_294_io_cout; // @[MUL.scala 102:19]
  wire  m_295_io_x1; // @[MUL.scala 102:19]
  wire  m_295_io_x2; // @[MUL.scala 102:19]
  wire  m_295_io_x3; // @[MUL.scala 102:19]
  wire  m_295_io_s; // @[MUL.scala 102:19]
  wire  m_295_io_cout; // @[MUL.scala 102:19]
  wire  m_296_io_x1; // @[MUL.scala 102:19]
  wire  m_296_io_x2; // @[MUL.scala 102:19]
  wire  m_296_io_x3; // @[MUL.scala 102:19]
  wire  m_296_io_s; // @[MUL.scala 102:19]
  wire  m_296_io_cout; // @[MUL.scala 102:19]
  wire  m_297_io_x1; // @[MUL.scala 102:19]
  wire  m_297_io_x2; // @[MUL.scala 102:19]
  wire  m_297_io_x3; // @[MUL.scala 102:19]
  wire  m_297_io_s; // @[MUL.scala 102:19]
  wire  m_297_io_cout; // @[MUL.scala 102:19]
  wire  m_298_io_x1; // @[MUL.scala 102:19]
  wire  m_298_io_x2; // @[MUL.scala 102:19]
  wire  m_298_io_x3; // @[MUL.scala 102:19]
  wire  m_298_io_s; // @[MUL.scala 102:19]
  wire  m_298_io_cout; // @[MUL.scala 102:19]
  wire  m_299_io_x1; // @[MUL.scala 102:19]
  wire  m_299_io_x2; // @[MUL.scala 102:19]
  wire  m_299_io_x3; // @[MUL.scala 102:19]
  wire  m_299_io_s; // @[MUL.scala 102:19]
  wire  m_299_io_cout; // @[MUL.scala 102:19]
  wire  m_300_io_x1; // @[MUL.scala 102:19]
  wire  m_300_io_x2; // @[MUL.scala 102:19]
  wire  m_300_io_x3; // @[MUL.scala 102:19]
  wire  m_300_io_s; // @[MUL.scala 102:19]
  wire  m_300_io_cout; // @[MUL.scala 102:19]
  wire  m_301_io_x1; // @[MUL.scala 102:19]
  wire  m_301_io_x2; // @[MUL.scala 102:19]
  wire  m_301_io_x3; // @[MUL.scala 102:19]
  wire  m_301_io_s; // @[MUL.scala 102:19]
  wire  m_301_io_cout; // @[MUL.scala 102:19]
  wire  m_302_io_x1; // @[MUL.scala 102:19]
  wire  m_302_io_x2; // @[MUL.scala 102:19]
  wire  m_302_io_x3; // @[MUL.scala 102:19]
  wire  m_302_io_s; // @[MUL.scala 102:19]
  wire  m_302_io_cout; // @[MUL.scala 102:19]
  wire  m_303_io_x1; // @[MUL.scala 102:19]
  wire  m_303_io_x2; // @[MUL.scala 102:19]
  wire  m_303_io_x3; // @[MUL.scala 102:19]
  wire  m_303_io_s; // @[MUL.scala 102:19]
  wire  m_303_io_cout; // @[MUL.scala 102:19]
  wire  m_304_io_x1; // @[MUL.scala 102:19]
  wire  m_304_io_x2; // @[MUL.scala 102:19]
  wire  m_304_io_x3; // @[MUL.scala 102:19]
  wire  m_304_io_s; // @[MUL.scala 102:19]
  wire  m_304_io_cout; // @[MUL.scala 102:19]
  wire  m_305_io_x1; // @[MUL.scala 102:19]
  wire  m_305_io_x2; // @[MUL.scala 102:19]
  wire  m_305_io_x3; // @[MUL.scala 102:19]
  wire  m_305_io_s; // @[MUL.scala 102:19]
  wire  m_305_io_cout; // @[MUL.scala 102:19]
  wire  m_306_io_x1; // @[MUL.scala 102:19]
  wire  m_306_io_x2; // @[MUL.scala 102:19]
  wire  m_306_io_x3; // @[MUL.scala 102:19]
  wire  m_306_io_s; // @[MUL.scala 102:19]
  wire  m_306_io_cout; // @[MUL.scala 102:19]
  wire  m_307_io_x1; // @[MUL.scala 102:19]
  wire  m_307_io_x2; // @[MUL.scala 102:19]
  wire  m_307_io_x3; // @[MUL.scala 102:19]
  wire  m_307_io_s; // @[MUL.scala 102:19]
  wire  m_307_io_cout; // @[MUL.scala 102:19]
  wire  m_308_io_x1; // @[MUL.scala 102:19]
  wire  m_308_io_x2; // @[MUL.scala 102:19]
  wire  m_308_io_x3; // @[MUL.scala 102:19]
  wire  m_308_io_s; // @[MUL.scala 102:19]
  wire  m_308_io_cout; // @[MUL.scala 102:19]
  wire  m_309_io_x1; // @[MUL.scala 102:19]
  wire  m_309_io_x2; // @[MUL.scala 102:19]
  wire  m_309_io_x3; // @[MUL.scala 102:19]
  wire  m_309_io_s; // @[MUL.scala 102:19]
  wire  m_309_io_cout; // @[MUL.scala 102:19]
  wire  m_310_io_x1; // @[MUL.scala 102:19]
  wire  m_310_io_x2; // @[MUL.scala 102:19]
  wire  m_310_io_x3; // @[MUL.scala 102:19]
  wire  m_310_io_s; // @[MUL.scala 102:19]
  wire  m_310_io_cout; // @[MUL.scala 102:19]
  wire  m_311_io_x1; // @[MUL.scala 102:19]
  wire  m_311_io_x2; // @[MUL.scala 102:19]
  wire  m_311_io_x3; // @[MUL.scala 102:19]
  wire  m_311_io_s; // @[MUL.scala 102:19]
  wire  m_311_io_cout; // @[MUL.scala 102:19]
  wire  m_312_io_in_0; // @[MUL.scala 124:19]
  wire  m_312_io_in_1; // @[MUL.scala 124:19]
  wire  m_312_io_out_0; // @[MUL.scala 124:19]
  wire  m_312_io_out_1; // @[MUL.scala 124:19]
  wire  m_313_io_x1; // @[MUL.scala 102:19]
  wire  m_313_io_x2; // @[MUL.scala 102:19]
  wire  m_313_io_x3; // @[MUL.scala 102:19]
  wire  m_313_io_s; // @[MUL.scala 102:19]
  wire  m_313_io_cout; // @[MUL.scala 102:19]
  wire  m_314_io_x1; // @[MUL.scala 102:19]
  wire  m_314_io_x2; // @[MUL.scala 102:19]
  wire  m_314_io_x3; // @[MUL.scala 102:19]
  wire  m_314_io_s; // @[MUL.scala 102:19]
  wire  m_314_io_cout; // @[MUL.scala 102:19]
  wire  m_315_io_x1; // @[MUL.scala 102:19]
  wire  m_315_io_x2; // @[MUL.scala 102:19]
  wire  m_315_io_x3; // @[MUL.scala 102:19]
  wire  m_315_io_s; // @[MUL.scala 102:19]
  wire  m_315_io_cout; // @[MUL.scala 102:19]
  wire  m_316_io_x1; // @[MUL.scala 102:19]
  wire  m_316_io_x2; // @[MUL.scala 102:19]
  wire  m_316_io_x3; // @[MUL.scala 102:19]
  wire  m_316_io_s; // @[MUL.scala 102:19]
  wire  m_316_io_cout; // @[MUL.scala 102:19]
  wire  m_317_io_x1; // @[MUL.scala 102:19]
  wire  m_317_io_x2; // @[MUL.scala 102:19]
  wire  m_317_io_x3; // @[MUL.scala 102:19]
  wire  m_317_io_s; // @[MUL.scala 102:19]
  wire  m_317_io_cout; // @[MUL.scala 102:19]
  wire  m_318_io_x1; // @[MUL.scala 102:19]
  wire  m_318_io_x2; // @[MUL.scala 102:19]
  wire  m_318_io_x3; // @[MUL.scala 102:19]
  wire  m_318_io_s; // @[MUL.scala 102:19]
  wire  m_318_io_cout; // @[MUL.scala 102:19]
  wire  m_319_io_x1; // @[MUL.scala 102:19]
  wire  m_319_io_x2; // @[MUL.scala 102:19]
  wire  m_319_io_x3; // @[MUL.scala 102:19]
  wire  m_319_io_s; // @[MUL.scala 102:19]
  wire  m_319_io_cout; // @[MUL.scala 102:19]
  wire  m_320_io_x1; // @[MUL.scala 102:19]
  wire  m_320_io_x2; // @[MUL.scala 102:19]
  wire  m_320_io_x3; // @[MUL.scala 102:19]
  wire  m_320_io_s; // @[MUL.scala 102:19]
  wire  m_320_io_cout; // @[MUL.scala 102:19]
  wire  m_321_io_x1; // @[MUL.scala 102:19]
  wire  m_321_io_x2; // @[MUL.scala 102:19]
  wire  m_321_io_x3; // @[MUL.scala 102:19]
  wire  m_321_io_s; // @[MUL.scala 102:19]
  wire  m_321_io_cout; // @[MUL.scala 102:19]
  wire  m_322_io_in_0; // @[MUL.scala 124:19]
  wire  m_322_io_in_1; // @[MUL.scala 124:19]
  wire  m_322_io_out_0; // @[MUL.scala 124:19]
  wire  m_322_io_out_1; // @[MUL.scala 124:19]
  wire  m_323_io_x1; // @[MUL.scala 102:19]
  wire  m_323_io_x2; // @[MUL.scala 102:19]
  wire  m_323_io_x3; // @[MUL.scala 102:19]
  wire  m_323_io_s; // @[MUL.scala 102:19]
  wire  m_323_io_cout; // @[MUL.scala 102:19]
  wire  m_324_io_x1; // @[MUL.scala 102:19]
  wire  m_324_io_x2; // @[MUL.scala 102:19]
  wire  m_324_io_x3; // @[MUL.scala 102:19]
  wire  m_324_io_s; // @[MUL.scala 102:19]
  wire  m_324_io_cout; // @[MUL.scala 102:19]
  wire  m_325_io_x1; // @[MUL.scala 102:19]
  wire  m_325_io_x2; // @[MUL.scala 102:19]
  wire  m_325_io_x3; // @[MUL.scala 102:19]
  wire  m_325_io_s; // @[MUL.scala 102:19]
  wire  m_325_io_cout; // @[MUL.scala 102:19]
  wire  m_326_io_x1; // @[MUL.scala 102:19]
  wire  m_326_io_x2; // @[MUL.scala 102:19]
  wire  m_326_io_x3; // @[MUL.scala 102:19]
  wire  m_326_io_s; // @[MUL.scala 102:19]
  wire  m_326_io_cout; // @[MUL.scala 102:19]
  wire  m_327_io_x1; // @[MUL.scala 102:19]
  wire  m_327_io_x2; // @[MUL.scala 102:19]
  wire  m_327_io_x3; // @[MUL.scala 102:19]
  wire  m_327_io_s; // @[MUL.scala 102:19]
  wire  m_327_io_cout; // @[MUL.scala 102:19]
  wire  m_328_io_x1; // @[MUL.scala 102:19]
  wire  m_328_io_x2; // @[MUL.scala 102:19]
  wire  m_328_io_x3; // @[MUL.scala 102:19]
  wire  m_328_io_s; // @[MUL.scala 102:19]
  wire  m_328_io_cout; // @[MUL.scala 102:19]
  wire  m_329_io_x1; // @[MUL.scala 102:19]
  wire  m_329_io_x2; // @[MUL.scala 102:19]
  wire  m_329_io_x3; // @[MUL.scala 102:19]
  wire  m_329_io_s; // @[MUL.scala 102:19]
  wire  m_329_io_cout; // @[MUL.scala 102:19]
  wire  m_330_io_x1; // @[MUL.scala 102:19]
  wire  m_330_io_x2; // @[MUL.scala 102:19]
  wire  m_330_io_x3; // @[MUL.scala 102:19]
  wire  m_330_io_s; // @[MUL.scala 102:19]
  wire  m_330_io_cout; // @[MUL.scala 102:19]
  wire  m_331_io_x1; // @[MUL.scala 102:19]
  wire  m_331_io_x2; // @[MUL.scala 102:19]
  wire  m_331_io_x3; // @[MUL.scala 102:19]
  wire  m_331_io_s; // @[MUL.scala 102:19]
  wire  m_331_io_cout; // @[MUL.scala 102:19]
  wire  m_332_io_x1; // @[MUL.scala 102:19]
  wire  m_332_io_x2; // @[MUL.scala 102:19]
  wire  m_332_io_x3; // @[MUL.scala 102:19]
  wire  m_332_io_s; // @[MUL.scala 102:19]
  wire  m_332_io_cout; // @[MUL.scala 102:19]
  wire  m_333_io_x1; // @[MUL.scala 102:19]
  wire  m_333_io_x2; // @[MUL.scala 102:19]
  wire  m_333_io_x3; // @[MUL.scala 102:19]
  wire  m_333_io_s; // @[MUL.scala 102:19]
  wire  m_333_io_cout; // @[MUL.scala 102:19]
  wire  m_334_io_x1; // @[MUL.scala 102:19]
  wire  m_334_io_x2; // @[MUL.scala 102:19]
  wire  m_334_io_x3; // @[MUL.scala 102:19]
  wire  m_334_io_s; // @[MUL.scala 102:19]
  wire  m_334_io_cout; // @[MUL.scala 102:19]
  wire  m_335_io_x1; // @[MUL.scala 102:19]
  wire  m_335_io_x2; // @[MUL.scala 102:19]
  wire  m_335_io_x3; // @[MUL.scala 102:19]
  wire  m_335_io_s; // @[MUL.scala 102:19]
  wire  m_335_io_cout; // @[MUL.scala 102:19]
  wire  m_336_io_x1; // @[MUL.scala 102:19]
  wire  m_336_io_x2; // @[MUL.scala 102:19]
  wire  m_336_io_x3; // @[MUL.scala 102:19]
  wire  m_336_io_s; // @[MUL.scala 102:19]
  wire  m_336_io_cout; // @[MUL.scala 102:19]
  wire  m_337_io_x1; // @[MUL.scala 102:19]
  wire  m_337_io_x2; // @[MUL.scala 102:19]
  wire  m_337_io_x3; // @[MUL.scala 102:19]
  wire  m_337_io_s; // @[MUL.scala 102:19]
  wire  m_337_io_cout; // @[MUL.scala 102:19]
  wire  m_338_io_x1; // @[MUL.scala 102:19]
  wire  m_338_io_x2; // @[MUL.scala 102:19]
  wire  m_338_io_x3; // @[MUL.scala 102:19]
  wire  m_338_io_s; // @[MUL.scala 102:19]
  wire  m_338_io_cout; // @[MUL.scala 102:19]
  wire  m_339_io_x1; // @[MUL.scala 102:19]
  wire  m_339_io_x2; // @[MUL.scala 102:19]
  wire  m_339_io_x3; // @[MUL.scala 102:19]
  wire  m_339_io_s; // @[MUL.scala 102:19]
  wire  m_339_io_cout; // @[MUL.scala 102:19]
  wire  m_340_io_x1; // @[MUL.scala 102:19]
  wire  m_340_io_x2; // @[MUL.scala 102:19]
  wire  m_340_io_x3; // @[MUL.scala 102:19]
  wire  m_340_io_s; // @[MUL.scala 102:19]
  wire  m_340_io_cout; // @[MUL.scala 102:19]
  wire  m_341_io_x1; // @[MUL.scala 102:19]
  wire  m_341_io_x2; // @[MUL.scala 102:19]
  wire  m_341_io_x3; // @[MUL.scala 102:19]
  wire  m_341_io_s; // @[MUL.scala 102:19]
  wire  m_341_io_cout; // @[MUL.scala 102:19]
  wire  m_342_io_x1; // @[MUL.scala 102:19]
  wire  m_342_io_x2; // @[MUL.scala 102:19]
  wire  m_342_io_x3; // @[MUL.scala 102:19]
  wire  m_342_io_s; // @[MUL.scala 102:19]
  wire  m_342_io_cout; // @[MUL.scala 102:19]
  wire  m_343_io_x1; // @[MUL.scala 102:19]
  wire  m_343_io_x2; // @[MUL.scala 102:19]
  wire  m_343_io_x3; // @[MUL.scala 102:19]
  wire  m_343_io_s; // @[MUL.scala 102:19]
  wire  m_343_io_cout; // @[MUL.scala 102:19]
  wire  m_344_io_x1; // @[MUL.scala 102:19]
  wire  m_344_io_x2; // @[MUL.scala 102:19]
  wire  m_344_io_x3; // @[MUL.scala 102:19]
  wire  m_344_io_s; // @[MUL.scala 102:19]
  wire  m_344_io_cout; // @[MUL.scala 102:19]
  wire  m_345_io_x1; // @[MUL.scala 102:19]
  wire  m_345_io_x2; // @[MUL.scala 102:19]
  wire  m_345_io_x3; // @[MUL.scala 102:19]
  wire  m_345_io_s; // @[MUL.scala 102:19]
  wire  m_345_io_cout; // @[MUL.scala 102:19]
  wire  m_346_io_x1; // @[MUL.scala 102:19]
  wire  m_346_io_x2; // @[MUL.scala 102:19]
  wire  m_346_io_x3; // @[MUL.scala 102:19]
  wire  m_346_io_s; // @[MUL.scala 102:19]
  wire  m_346_io_cout; // @[MUL.scala 102:19]
  wire  m_347_io_x1; // @[MUL.scala 102:19]
  wire  m_347_io_x2; // @[MUL.scala 102:19]
  wire  m_347_io_x3; // @[MUL.scala 102:19]
  wire  m_347_io_s; // @[MUL.scala 102:19]
  wire  m_347_io_cout; // @[MUL.scala 102:19]
  wire  m_348_io_x1; // @[MUL.scala 102:19]
  wire  m_348_io_x2; // @[MUL.scala 102:19]
  wire  m_348_io_x3; // @[MUL.scala 102:19]
  wire  m_348_io_s; // @[MUL.scala 102:19]
  wire  m_348_io_cout; // @[MUL.scala 102:19]
  wire  m_349_io_x1; // @[MUL.scala 102:19]
  wire  m_349_io_x2; // @[MUL.scala 102:19]
  wire  m_349_io_x3; // @[MUL.scala 102:19]
  wire  m_349_io_s; // @[MUL.scala 102:19]
  wire  m_349_io_cout; // @[MUL.scala 102:19]
  wire  m_350_io_x1; // @[MUL.scala 102:19]
  wire  m_350_io_x2; // @[MUL.scala 102:19]
  wire  m_350_io_x3; // @[MUL.scala 102:19]
  wire  m_350_io_s; // @[MUL.scala 102:19]
  wire  m_350_io_cout; // @[MUL.scala 102:19]
  wire  m_351_io_x1; // @[MUL.scala 102:19]
  wire  m_351_io_x2; // @[MUL.scala 102:19]
  wire  m_351_io_x3; // @[MUL.scala 102:19]
  wire  m_351_io_s; // @[MUL.scala 102:19]
  wire  m_351_io_cout; // @[MUL.scala 102:19]
  wire  m_352_io_x1; // @[MUL.scala 102:19]
  wire  m_352_io_x2; // @[MUL.scala 102:19]
  wire  m_352_io_x3; // @[MUL.scala 102:19]
  wire  m_352_io_s; // @[MUL.scala 102:19]
  wire  m_352_io_cout; // @[MUL.scala 102:19]
  wire  m_353_io_x1; // @[MUL.scala 102:19]
  wire  m_353_io_x2; // @[MUL.scala 102:19]
  wire  m_353_io_x3; // @[MUL.scala 102:19]
  wire  m_353_io_s; // @[MUL.scala 102:19]
  wire  m_353_io_cout; // @[MUL.scala 102:19]
  wire  m_354_io_x1; // @[MUL.scala 102:19]
  wire  m_354_io_x2; // @[MUL.scala 102:19]
  wire  m_354_io_x3; // @[MUL.scala 102:19]
  wire  m_354_io_s; // @[MUL.scala 102:19]
  wire  m_354_io_cout; // @[MUL.scala 102:19]
  wire  m_355_io_x1; // @[MUL.scala 102:19]
  wire  m_355_io_x2; // @[MUL.scala 102:19]
  wire  m_355_io_x3; // @[MUL.scala 102:19]
  wire  m_355_io_s; // @[MUL.scala 102:19]
  wire  m_355_io_cout; // @[MUL.scala 102:19]
  wire  m_356_io_x1; // @[MUL.scala 102:19]
  wire  m_356_io_x2; // @[MUL.scala 102:19]
  wire  m_356_io_x3; // @[MUL.scala 102:19]
  wire  m_356_io_s; // @[MUL.scala 102:19]
  wire  m_356_io_cout; // @[MUL.scala 102:19]
  wire  m_357_io_x1; // @[MUL.scala 102:19]
  wire  m_357_io_x2; // @[MUL.scala 102:19]
  wire  m_357_io_x3; // @[MUL.scala 102:19]
  wire  m_357_io_s; // @[MUL.scala 102:19]
  wire  m_357_io_cout; // @[MUL.scala 102:19]
  wire  m_358_io_x1; // @[MUL.scala 102:19]
  wire  m_358_io_x2; // @[MUL.scala 102:19]
  wire  m_358_io_x3; // @[MUL.scala 102:19]
  wire  m_358_io_s; // @[MUL.scala 102:19]
  wire  m_358_io_cout; // @[MUL.scala 102:19]
  wire  m_359_io_x1; // @[MUL.scala 102:19]
  wire  m_359_io_x2; // @[MUL.scala 102:19]
  wire  m_359_io_x3; // @[MUL.scala 102:19]
  wire  m_359_io_s; // @[MUL.scala 102:19]
  wire  m_359_io_cout; // @[MUL.scala 102:19]
  wire  m_360_io_x1; // @[MUL.scala 102:19]
  wire  m_360_io_x2; // @[MUL.scala 102:19]
  wire  m_360_io_x3; // @[MUL.scala 102:19]
  wire  m_360_io_s; // @[MUL.scala 102:19]
  wire  m_360_io_cout; // @[MUL.scala 102:19]
  wire  m_361_io_x1; // @[MUL.scala 102:19]
  wire  m_361_io_x2; // @[MUL.scala 102:19]
  wire  m_361_io_x3; // @[MUL.scala 102:19]
  wire  m_361_io_s; // @[MUL.scala 102:19]
  wire  m_361_io_cout; // @[MUL.scala 102:19]
  wire  m_362_io_x1; // @[MUL.scala 102:19]
  wire  m_362_io_x2; // @[MUL.scala 102:19]
  wire  m_362_io_x3; // @[MUL.scala 102:19]
  wire  m_362_io_s; // @[MUL.scala 102:19]
  wire  m_362_io_cout; // @[MUL.scala 102:19]
  wire  m_363_io_x1; // @[MUL.scala 102:19]
  wire  m_363_io_x2; // @[MUL.scala 102:19]
  wire  m_363_io_x3; // @[MUL.scala 102:19]
  wire  m_363_io_s; // @[MUL.scala 102:19]
  wire  m_363_io_cout; // @[MUL.scala 102:19]
  wire  m_364_io_x1; // @[MUL.scala 102:19]
  wire  m_364_io_x2; // @[MUL.scala 102:19]
  wire  m_364_io_x3; // @[MUL.scala 102:19]
  wire  m_364_io_s; // @[MUL.scala 102:19]
  wire  m_364_io_cout; // @[MUL.scala 102:19]
  wire  m_365_io_x1; // @[MUL.scala 102:19]
  wire  m_365_io_x2; // @[MUL.scala 102:19]
  wire  m_365_io_x3; // @[MUL.scala 102:19]
  wire  m_365_io_s; // @[MUL.scala 102:19]
  wire  m_365_io_cout; // @[MUL.scala 102:19]
  wire  m_366_io_x1; // @[MUL.scala 102:19]
  wire  m_366_io_x2; // @[MUL.scala 102:19]
  wire  m_366_io_x3; // @[MUL.scala 102:19]
  wire  m_366_io_s; // @[MUL.scala 102:19]
  wire  m_366_io_cout; // @[MUL.scala 102:19]
  wire  m_367_io_x1; // @[MUL.scala 102:19]
  wire  m_367_io_x2; // @[MUL.scala 102:19]
  wire  m_367_io_x3; // @[MUL.scala 102:19]
  wire  m_367_io_s; // @[MUL.scala 102:19]
  wire  m_367_io_cout; // @[MUL.scala 102:19]
  wire  m_368_io_x1; // @[MUL.scala 102:19]
  wire  m_368_io_x2; // @[MUL.scala 102:19]
  wire  m_368_io_x3; // @[MUL.scala 102:19]
  wire  m_368_io_s; // @[MUL.scala 102:19]
  wire  m_368_io_cout; // @[MUL.scala 102:19]
  wire  m_369_io_x1; // @[MUL.scala 102:19]
  wire  m_369_io_x2; // @[MUL.scala 102:19]
  wire  m_369_io_x3; // @[MUL.scala 102:19]
  wire  m_369_io_s; // @[MUL.scala 102:19]
  wire  m_369_io_cout; // @[MUL.scala 102:19]
  wire  m_370_io_x1; // @[MUL.scala 102:19]
  wire  m_370_io_x2; // @[MUL.scala 102:19]
  wire  m_370_io_x3; // @[MUL.scala 102:19]
  wire  m_370_io_s; // @[MUL.scala 102:19]
  wire  m_370_io_cout; // @[MUL.scala 102:19]
  wire  m_371_io_x1; // @[MUL.scala 102:19]
  wire  m_371_io_x2; // @[MUL.scala 102:19]
  wire  m_371_io_x3; // @[MUL.scala 102:19]
  wire  m_371_io_s; // @[MUL.scala 102:19]
  wire  m_371_io_cout; // @[MUL.scala 102:19]
  wire  m_372_io_x1; // @[MUL.scala 102:19]
  wire  m_372_io_x2; // @[MUL.scala 102:19]
  wire  m_372_io_x3; // @[MUL.scala 102:19]
  wire  m_372_io_s; // @[MUL.scala 102:19]
  wire  m_372_io_cout; // @[MUL.scala 102:19]
  wire  m_373_io_in_0; // @[MUL.scala 124:19]
  wire  m_373_io_in_1; // @[MUL.scala 124:19]
  wire  m_373_io_out_0; // @[MUL.scala 124:19]
  wire  m_373_io_out_1; // @[MUL.scala 124:19]
  wire  m_374_io_x1; // @[MUL.scala 102:19]
  wire  m_374_io_x2; // @[MUL.scala 102:19]
  wire  m_374_io_x3; // @[MUL.scala 102:19]
  wire  m_374_io_s; // @[MUL.scala 102:19]
  wire  m_374_io_cout; // @[MUL.scala 102:19]
  wire  m_375_io_x1; // @[MUL.scala 102:19]
  wire  m_375_io_x2; // @[MUL.scala 102:19]
  wire  m_375_io_x3; // @[MUL.scala 102:19]
  wire  m_375_io_s; // @[MUL.scala 102:19]
  wire  m_375_io_cout; // @[MUL.scala 102:19]
  wire  m_376_io_x1; // @[MUL.scala 102:19]
  wire  m_376_io_x2; // @[MUL.scala 102:19]
  wire  m_376_io_x3; // @[MUL.scala 102:19]
  wire  m_376_io_s; // @[MUL.scala 102:19]
  wire  m_376_io_cout; // @[MUL.scala 102:19]
  wire  m_377_io_x1; // @[MUL.scala 102:19]
  wire  m_377_io_x2; // @[MUL.scala 102:19]
  wire  m_377_io_x3; // @[MUL.scala 102:19]
  wire  m_377_io_s; // @[MUL.scala 102:19]
  wire  m_377_io_cout; // @[MUL.scala 102:19]
  wire  m_378_io_x1; // @[MUL.scala 102:19]
  wire  m_378_io_x2; // @[MUL.scala 102:19]
  wire  m_378_io_x3; // @[MUL.scala 102:19]
  wire  m_378_io_s; // @[MUL.scala 102:19]
  wire  m_378_io_cout; // @[MUL.scala 102:19]
  wire  m_379_io_x1; // @[MUL.scala 102:19]
  wire  m_379_io_x2; // @[MUL.scala 102:19]
  wire  m_379_io_x3; // @[MUL.scala 102:19]
  wire  m_379_io_s; // @[MUL.scala 102:19]
  wire  m_379_io_cout; // @[MUL.scala 102:19]
  wire  m_380_io_x1; // @[MUL.scala 102:19]
  wire  m_380_io_x2; // @[MUL.scala 102:19]
  wire  m_380_io_x3; // @[MUL.scala 102:19]
  wire  m_380_io_s; // @[MUL.scala 102:19]
  wire  m_380_io_cout; // @[MUL.scala 102:19]
  wire  m_381_io_x1; // @[MUL.scala 102:19]
  wire  m_381_io_x2; // @[MUL.scala 102:19]
  wire  m_381_io_x3; // @[MUL.scala 102:19]
  wire  m_381_io_s; // @[MUL.scala 102:19]
  wire  m_381_io_cout; // @[MUL.scala 102:19]
  wire  m_382_io_x1; // @[MUL.scala 102:19]
  wire  m_382_io_x2; // @[MUL.scala 102:19]
  wire  m_382_io_x3; // @[MUL.scala 102:19]
  wire  m_382_io_s; // @[MUL.scala 102:19]
  wire  m_382_io_cout; // @[MUL.scala 102:19]
  wire  m_383_io_x1; // @[MUL.scala 102:19]
  wire  m_383_io_x2; // @[MUL.scala 102:19]
  wire  m_383_io_x3; // @[MUL.scala 102:19]
  wire  m_383_io_s; // @[MUL.scala 102:19]
  wire  m_383_io_cout; // @[MUL.scala 102:19]
  wire  m_384_io_in_0; // @[MUL.scala 124:19]
  wire  m_384_io_in_1; // @[MUL.scala 124:19]
  wire  m_384_io_out_0; // @[MUL.scala 124:19]
  wire  m_384_io_out_1; // @[MUL.scala 124:19]
  wire  m_385_io_x1; // @[MUL.scala 102:19]
  wire  m_385_io_x2; // @[MUL.scala 102:19]
  wire  m_385_io_x3; // @[MUL.scala 102:19]
  wire  m_385_io_s; // @[MUL.scala 102:19]
  wire  m_385_io_cout; // @[MUL.scala 102:19]
  wire  m_386_io_x1; // @[MUL.scala 102:19]
  wire  m_386_io_x2; // @[MUL.scala 102:19]
  wire  m_386_io_x3; // @[MUL.scala 102:19]
  wire  m_386_io_s; // @[MUL.scala 102:19]
  wire  m_386_io_cout; // @[MUL.scala 102:19]
  wire  m_387_io_x1; // @[MUL.scala 102:19]
  wire  m_387_io_x2; // @[MUL.scala 102:19]
  wire  m_387_io_x3; // @[MUL.scala 102:19]
  wire  m_387_io_s; // @[MUL.scala 102:19]
  wire  m_387_io_cout; // @[MUL.scala 102:19]
  wire  m_388_io_x1; // @[MUL.scala 102:19]
  wire  m_388_io_x2; // @[MUL.scala 102:19]
  wire  m_388_io_x3; // @[MUL.scala 102:19]
  wire  m_388_io_s; // @[MUL.scala 102:19]
  wire  m_388_io_cout; // @[MUL.scala 102:19]
  wire  m_389_io_x1; // @[MUL.scala 102:19]
  wire  m_389_io_x2; // @[MUL.scala 102:19]
  wire  m_389_io_x3; // @[MUL.scala 102:19]
  wire  m_389_io_s; // @[MUL.scala 102:19]
  wire  m_389_io_cout; // @[MUL.scala 102:19]
  wire  m_390_io_x1; // @[MUL.scala 102:19]
  wire  m_390_io_x2; // @[MUL.scala 102:19]
  wire  m_390_io_x3; // @[MUL.scala 102:19]
  wire  m_390_io_s; // @[MUL.scala 102:19]
  wire  m_390_io_cout; // @[MUL.scala 102:19]
  wire  m_391_io_x1; // @[MUL.scala 102:19]
  wire  m_391_io_x2; // @[MUL.scala 102:19]
  wire  m_391_io_x3; // @[MUL.scala 102:19]
  wire  m_391_io_s; // @[MUL.scala 102:19]
  wire  m_391_io_cout; // @[MUL.scala 102:19]
  wire  m_392_io_x1; // @[MUL.scala 102:19]
  wire  m_392_io_x2; // @[MUL.scala 102:19]
  wire  m_392_io_x3; // @[MUL.scala 102:19]
  wire  m_392_io_s; // @[MUL.scala 102:19]
  wire  m_392_io_cout; // @[MUL.scala 102:19]
  wire  m_393_io_x1; // @[MUL.scala 102:19]
  wire  m_393_io_x2; // @[MUL.scala 102:19]
  wire  m_393_io_x3; // @[MUL.scala 102:19]
  wire  m_393_io_s; // @[MUL.scala 102:19]
  wire  m_393_io_cout; // @[MUL.scala 102:19]
  wire  m_394_io_x1; // @[MUL.scala 102:19]
  wire  m_394_io_x2; // @[MUL.scala 102:19]
  wire  m_394_io_x3; // @[MUL.scala 102:19]
  wire  m_394_io_s; // @[MUL.scala 102:19]
  wire  m_394_io_cout; // @[MUL.scala 102:19]
  wire  m_395_io_x1; // @[MUL.scala 102:19]
  wire  m_395_io_x2; // @[MUL.scala 102:19]
  wire  m_395_io_x3; // @[MUL.scala 102:19]
  wire  m_395_io_s; // @[MUL.scala 102:19]
  wire  m_395_io_cout; // @[MUL.scala 102:19]
  wire  m_396_io_x1; // @[MUL.scala 102:19]
  wire  m_396_io_x2; // @[MUL.scala 102:19]
  wire  m_396_io_x3; // @[MUL.scala 102:19]
  wire  m_396_io_s; // @[MUL.scala 102:19]
  wire  m_396_io_cout; // @[MUL.scala 102:19]
  wire  m_397_io_x1; // @[MUL.scala 102:19]
  wire  m_397_io_x2; // @[MUL.scala 102:19]
  wire  m_397_io_x3; // @[MUL.scala 102:19]
  wire  m_397_io_s; // @[MUL.scala 102:19]
  wire  m_397_io_cout; // @[MUL.scala 102:19]
  wire  m_398_io_x1; // @[MUL.scala 102:19]
  wire  m_398_io_x2; // @[MUL.scala 102:19]
  wire  m_398_io_x3; // @[MUL.scala 102:19]
  wire  m_398_io_s; // @[MUL.scala 102:19]
  wire  m_398_io_cout; // @[MUL.scala 102:19]
  wire  m_399_io_x1; // @[MUL.scala 102:19]
  wire  m_399_io_x2; // @[MUL.scala 102:19]
  wire  m_399_io_x3; // @[MUL.scala 102:19]
  wire  m_399_io_s; // @[MUL.scala 102:19]
  wire  m_399_io_cout; // @[MUL.scala 102:19]
  wire  m_400_io_x1; // @[MUL.scala 102:19]
  wire  m_400_io_x2; // @[MUL.scala 102:19]
  wire  m_400_io_x3; // @[MUL.scala 102:19]
  wire  m_400_io_s; // @[MUL.scala 102:19]
  wire  m_400_io_cout; // @[MUL.scala 102:19]
  wire  m_401_io_x1; // @[MUL.scala 102:19]
  wire  m_401_io_x2; // @[MUL.scala 102:19]
  wire  m_401_io_x3; // @[MUL.scala 102:19]
  wire  m_401_io_s; // @[MUL.scala 102:19]
  wire  m_401_io_cout; // @[MUL.scala 102:19]
  wire  m_402_io_x1; // @[MUL.scala 102:19]
  wire  m_402_io_x2; // @[MUL.scala 102:19]
  wire  m_402_io_x3; // @[MUL.scala 102:19]
  wire  m_402_io_s; // @[MUL.scala 102:19]
  wire  m_402_io_cout; // @[MUL.scala 102:19]
  wire  m_403_io_x1; // @[MUL.scala 102:19]
  wire  m_403_io_x2; // @[MUL.scala 102:19]
  wire  m_403_io_x3; // @[MUL.scala 102:19]
  wire  m_403_io_s; // @[MUL.scala 102:19]
  wire  m_403_io_cout; // @[MUL.scala 102:19]
  wire  m_404_io_x1; // @[MUL.scala 102:19]
  wire  m_404_io_x2; // @[MUL.scala 102:19]
  wire  m_404_io_x3; // @[MUL.scala 102:19]
  wire  m_404_io_s; // @[MUL.scala 102:19]
  wire  m_404_io_cout; // @[MUL.scala 102:19]
  wire  m_405_io_x1; // @[MUL.scala 102:19]
  wire  m_405_io_x2; // @[MUL.scala 102:19]
  wire  m_405_io_x3; // @[MUL.scala 102:19]
  wire  m_405_io_s; // @[MUL.scala 102:19]
  wire  m_405_io_cout; // @[MUL.scala 102:19]
  wire  m_406_io_x1; // @[MUL.scala 102:19]
  wire  m_406_io_x2; // @[MUL.scala 102:19]
  wire  m_406_io_x3; // @[MUL.scala 102:19]
  wire  m_406_io_s; // @[MUL.scala 102:19]
  wire  m_406_io_cout; // @[MUL.scala 102:19]
  wire  m_407_io_x1; // @[MUL.scala 102:19]
  wire  m_407_io_x2; // @[MUL.scala 102:19]
  wire  m_407_io_x3; // @[MUL.scala 102:19]
  wire  m_407_io_s; // @[MUL.scala 102:19]
  wire  m_407_io_cout; // @[MUL.scala 102:19]
  wire  m_408_io_x1; // @[MUL.scala 102:19]
  wire  m_408_io_x2; // @[MUL.scala 102:19]
  wire  m_408_io_x3; // @[MUL.scala 102:19]
  wire  m_408_io_s; // @[MUL.scala 102:19]
  wire  m_408_io_cout; // @[MUL.scala 102:19]
  wire  m_409_io_x1; // @[MUL.scala 102:19]
  wire  m_409_io_x2; // @[MUL.scala 102:19]
  wire  m_409_io_x3; // @[MUL.scala 102:19]
  wire  m_409_io_s; // @[MUL.scala 102:19]
  wire  m_409_io_cout; // @[MUL.scala 102:19]
  wire  m_410_io_x1; // @[MUL.scala 102:19]
  wire  m_410_io_x2; // @[MUL.scala 102:19]
  wire  m_410_io_x3; // @[MUL.scala 102:19]
  wire  m_410_io_s; // @[MUL.scala 102:19]
  wire  m_410_io_cout; // @[MUL.scala 102:19]
  wire  m_411_io_x1; // @[MUL.scala 102:19]
  wire  m_411_io_x2; // @[MUL.scala 102:19]
  wire  m_411_io_x3; // @[MUL.scala 102:19]
  wire  m_411_io_s; // @[MUL.scala 102:19]
  wire  m_411_io_cout; // @[MUL.scala 102:19]
  wire  m_412_io_x1; // @[MUL.scala 102:19]
  wire  m_412_io_x2; // @[MUL.scala 102:19]
  wire  m_412_io_x3; // @[MUL.scala 102:19]
  wire  m_412_io_s; // @[MUL.scala 102:19]
  wire  m_412_io_cout; // @[MUL.scala 102:19]
  wire  m_413_io_x1; // @[MUL.scala 102:19]
  wire  m_413_io_x2; // @[MUL.scala 102:19]
  wire  m_413_io_x3; // @[MUL.scala 102:19]
  wire  m_413_io_s; // @[MUL.scala 102:19]
  wire  m_413_io_cout; // @[MUL.scala 102:19]
  wire  m_414_io_x1; // @[MUL.scala 102:19]
  wire  m_414_io_x2; // @[MUL.scala 102:19]
  wire  m_414_io_x3; // @[MUL.scala 102:19]
  wire  m_414_io_s; // @[MUL.scala 102:19]
  wire  m_414_io_cout; // @[MUL.scala 102:19]
  wire  m_415_io_x1; // @[MUL.scala 102:19]
  wire  m_415_io_x2; // @[MUL.scala 102:19]
  wire  m_415_io_x3; // @[MUL.scala 102:19]
  wire  m_415_io_s; // @[MUL.scala 102:19]
  wire  m_415_io_cout; // @[MUL.scala 102:19]
  wire  m_416_io_x1; // @[MUL.scala 102:19]
  wire  m_416_io_x2; // @[MUL.scala 102:19]
  wire  m_416_io_x3; // @[MUL.scala 102:19]
  wire  m_416_io_s; // @[MUL.scala 102:19]
  wire  m_416_io_cout; // @[MUL.scala 102:19]
  wire  m_417_io_x1; // @[MUL.scala 102:19]
  wire  m_417_io_x2; // @[MUL.scala 102:19]
  wire  m_417_io_x3; // @[MUL.scala 102:19]
  wire  m_417_io_s; // @[MUL.scala 102:19]
  wire  m_417_io_cout; // @[MUL.scala 102:19]
  wire  m_418_io_x1; // @[MUL.scala 102:19]
  wire  m_418_io_x2; // @[MUL.scala 102:19]
  wire  m_418_io_x3; // @[MUL.scala 102:19]
  wire  m_418_io_s; // @[MUL.scala 102:19]
  wire  m_418_io_cout; // @[MUL.scala 102:19]
  wire  m_419_io_x1; // @[MUL.scala 102:19]
  wire  m_419_io_x2; // @[MUL.scala 102:19]
  wire  m_419_io_x3; // @[MUL.scala 102:19]
  wire  m_419_io_s; // @[MUL.scala 102:19]
  wire  m_419_io_cout; // @[MUL.scala 102:19]
  wire  m_420_io_x1; // @[MUL.scala 102:19]
  wire  m_420_io_x2; // @[MUL.scala 102:19]
  wire  m_420_io_x3; // @[MUL.scala 102:19]
  wire  m_420_io_s; // @[MUL.scala 102:19]
  wire  m_420_io_cout; // @[MUL.scala 102:19]
  wire  m_421_io_x1; // @[MUL.scala 102:19]
  wire  m_421_io_x2; // @[MUL.scala 102:19]
  wire  m_421_io_x3; // @[MUL.scala 102:19]
  wire  m_421_io_s; // @[MUL.scala 102:19]
  wire  m_421_io_cout; // @[MUL.scala 102:19]
  wire  m_422_io_x1; // @[MUL.scala 102:19]
  wire  m_422_io_x2; // @[MUL.scala 102:19]
  wire  m_422_io_x3; // @[MUL.scala 102:19]
  wire  m_422_io_s; // @[MUL.scala 102:19]
  wire  m_422_io_cout; // @[MUL.scala 102:19]
  wire  m_423_io_x1; // @[MUL.scala 102:19]
  wire  m_423_io_x2; // @[MUL.scala 102:19]
  wire  m_423_io_x3; // @[MUL.scala 102:19]
  wire  m_423_io_s; // @[MUL.scala 102:19]
  wire  m_423_io_cout; // @[MUL.scala 102:19]
  wire  m_424_io_x1; // @[MUL.scala 102:19]
  wire  m_424_io_x2; // @[MUL.scala 102:19]
  wire  m_424_io_x3; // @[MUL.scala 102:19]
  wire  m_424_io_s; // @[MUL.scala 102:19]
  wire  m_424_io_cout; // @[MUL.scala 102:19]
  wire  m_425_io_x1; // @[MUL.scala 102:19]
  wire  m_425_io_x2; // @[MUL.scala 102:19]
  wire  m_425_io_x3; // @[MUL.scala 102:19]
  wire  m_425_io_s; // @[MUL.scala 102:19]
  wire  m_425_io_cout; // @[MUL.scala 102:19]
  wire  m_426_io_x1; // @[MUL.scala 102:19]
  wire  m_426_io_x2; // @[MUL.scala 102:19]
  wire  m_426_io_x3; // @[MUL.scala 102:19]
  wire  m_426_io_s; // @[MUL.scala 102:19]
  wire  m_426_io_cout; // @[MUL.scala 102:19]
  wire  m_427_io_x1; // @[MUL.scala 102:19]
  wire  m_427_io_x2; // @[MUL.scala 102:19]
  wire  m_427_io_x3; // @[MUL.scala 102:19]
  wire  m_427_io_s; // @[MUL.scala 102:19]
  wire  m_427_io_cout; // @[MUL.scala 102:19]
  wire  m_428_io_x1; // @[MUL.scala 102:19]
  wire  m_428_io_x2; // @[MUL.scala 102:19]
  wire  m_428_io_x3; // @[MUL.scala 102:19]
  wire  m_428_io_s; // @[MUL.scala 102:19]
  wire  m_428_io_cout; // @[MUL.scala 102:19]
  wire  m_429_io_x1; // @[MUL.scala 102:19]
  wire  m_429_io_x2; // @[MUL.scala 102:19]
  wire  m_429_io_x3; // @[MUL.scala 102:19]
  wire  m_429_io_s; // @[MUL.scala 102:19]
  wire  m_429_io_cout; // @[MUL.scala 102:19]
  wire  m_430_io_x1; // @[MUL.scala 102:19]
  wire  m_430_io_x2; // @[MUL.scala 102:19]
  wire  m_430_io_x3; // @[MUL.scala 102:19]
  wire  m_430_io_s; // @[MUL.scala 102:19]
  wire  m_430_io_cout; // @[MUL.scala 102:19]
  wire  m_431_io_x1; // @[MUL.scala 102:19]
  wire  m_431_io_x2; // @[MUL.scala 102:19]
  wire  m_431_io_x3; // @[MUL.scala 102:19]
  wire  m_431_io_s; // @[MUL.scala 102:19]
  wire  m_431_io_cout; // @[MUL.scala 102:19]
  wire  m_432_io_x1; // @[MUL.scala 102:19]
  wire  m_432_io_x2; // @[MUL.scala 102:19]
  wire  m_432_io_x3; // @[MUL.scala 102:19]
  wire  m_432_io_s; // @[MUL.scala 102:19]
  wire  m_432_io_cout; // @[MUL.scala 102:19]
  wire  m_433_io_x1; // @[MUL.scala 102:19]
  wire  m_433_io_x2; // @[MUL.scala 102:19]
  wire  m_433_io_x3; // @[MUL.scala 102:19]
  wire  m_433_io_s; // @[MUL.scala 102:19]
  wire  m_433_io_cout; // @[MUL.scala 102:19]
  wire  m_434_io_x1; // @[MUL.scala 102:19]
  wire  m_434_io_x2; // @[MUL.scala 102:19]
  wire  m_434_io_x3; // @[MUL.scala 102:19]
  wire  m_434_io_s; // @[MUL.scala 102:19]
  wire  m_434_io_cout; // @[MUL.scala 102:19]
  wire  m_435_io_x1; // @[MUL.scala 102:19]
  wire  m_435_io_x2; // @[MUL.scala 102:19]
  wire  m_435_io_x3; // @[MUL.scala 102:19]
  wire  m_435_io_s; // @[MUL.scala 102:19]
  wire  m_435_io_cout; // @[MUL.scala 102:19]
  wire  m_436_io_x1; // @[MUL.scala 102:19]
  wire  m_436_io_x2; // @[MUL.scala 102:19]
  wire  m_436_io_x3; // @[MUL.scala 102:19]
  wire  m_436_io_s; // @[MUL.scala 102:19]
  wire  m_436_io_cout; // @[MUL.scala 102:19]
  wire  m_437_io_x1; // @[MUL.scala 102:19]
  wire  m_437_io_x2; // @[MUL.scala 102:19]
  wire  m_437_io_x3; // @[MUL.scala 102:19]
  wire  m_437_io_s; // @[MUL.scala 102:19]
  wire  m_437_io_cout; // @[MUL.scala 102:19]
  wire  m_438_io_x1; // @[MUL.scala 102:19]
  wire  m_438_io_x2; // @[MUL.scala 102:19]
  wire  m_438_io_x3; // @[MUL.scala 102:19]
  wire  m_438_io_s; // @[MUL.scala 102:19]
  wire  m_438_io_cout; // @[MUL.scala 102:19]
  wire  m_439_io_x1; // @[MUL.scala 102:19]
  wire  m_439_io_x2; // @[MUL.scala 102:19]
  wire  m_439_io_x3; // @[MUL.scala 102:19]
  wire  m_439_io_s; // @[MUL.scala 102:19]
  wire  m_439_io_cout; // @[MUL.scala 102:19]
  wire  m_440_io_x1; // @[MUL.scala 102:19]
  wire  m_440_io_x2; // @[MUL.scala 102:19]
  wire  m_440_io_x3; // @[MUL.scala 102:19]
  wire  m_440_io_s; // @[MUL.scala 102:19]
  wire  m_440_io_cout; // @[MUL.scala 102:19]
  wire  m_441_io_x1; // @[MUL.scala 102:19]
  wire  m_441_io_x2; // @[MUL.scala 102:19]
  wire  m_441_io_x3; // @[MUL.scala 102:19]
  wire  m_441_io_s; // @[MUL.scala 102:19]
  wire  m_441_io_cout; // @[MUL.scala 102:19]
  wire  m_442_io_x1; // @[MUL.scala 102:19]
  wire  m_442_io_x2; // @[MUL.scala 102:19]
  wire  m_442_io_x3; // @[MUL.scala 102:19]
  wire  m_442_io_s; // @[MUL.scala 102:19]
  wire  m_442_io_cout; // @[MUL.scala 102:19]
  wire  m_443_io_x1; // @[MUL.scala 102:19]
  wire  m_443_io_x2; // @[MUL.scala 102:19]
  wire  m_443_io_x3; // @[MUL.scala 102:19]
  wire  m_443_io_s; // @[MUL.scala 102:19]
  wire  m_443_io_cout; // @[MUL.scala 102:19]
  wire  m_444_io_x1; // @[MUL.scala 102:19]
  wire  m_444_io_x2; // @[MUL.scala 102:19]
  wire  m_444_io_x3; // @[MUL.scala 102:19]
  wire  m_444_io_s; // @[MUL.scala 102:19]
  wire  m_444_io_cout; // @[MUL.scala 102:19]
  wire  m_445_io_x1; // @[MUL.scala 102:19]
  wire  m_445_io_x2; // @[MUL.scala 102:19]
  wire  m_445_io_x3; // @[MUL.scala 102:19]
  wire  m_445_io_s; // @[MUL.scala 102:19]
  wire  m_445_io_cout; // @[MUL.scala 102:19]
  wire  m_446_io_x1; // @[MUL.scala 102:19]
  wire  m_446_io_x2; // @[MUL.scala 102:19]
  wire  m_446_io_x3; // @[MUL.scala 102:19]
  wire  m_446_io_s; // @[MUL.scala 102:19]
  wire  m_446_io_cout; // @[MUL.scala 102:19]
  wire  m_447_io_x1; // @[MUL.scala 102:19]
  wire  m_447_io_x2; // @[MUL.scala 102:19]
  wire  m_447_io_x3; // @[MUL.scala 102:19]
  wire  m_447_io_s; // @[MUL.scala 102:19]
  wire  m_447_io_cout; // @[MUL.scala 102:19]
  wire  m_448_io_x1; // @[MUL.scala 102:19]
  wire  m_448_io_x2; // @[MUL.scala 102:19]
  wire  m_448_io_x3; // @[MUL.scala 102:19]
  wire  m_448_io_s; // @[MUL.scala 102:19]
  wire  m_448_io_cout; // @[MUL.scala 102:19]
  wire  m_449_io_x1; // @[MUL.scala 102:19]
  wire  m_449_io_x2; // @[MUL.scala 102:19]
  wire  m_449_io_x3; // @[MUL.scala 102:19]
  wire  m_449_io_s; // @[MUL.scala 102:19]
  wire  m_449_io_cout; // @[MUL.scala 102:19]
  wire  m_450_io_x1; // @[MUL.scala 102:19]
  wire  m_450_io_x2; // @[MUL.scala 102:19]
  wire  m_450_io_x3; // @[MUL.scala 102:19]
  wire  m_450_io_s; // @[MUL.scala 102:19]
  wire  m_450_io_cout; // @[MUL.scala 102:19]
  wire  m_451_io_x1; // @[MUL.scala 102:19]
  wire  m_451_io_x2; // @[MUL.scala 102:19]
  wire  m_451_io_x3; // @[MUL.scala 102:19]
  wire  m_451_io_s; // @[MUL.scala 102:19]
  wire  m_451_io_cout; // @[MUL.scala 102:19]
  wire  m_452_io_x1; // @[MUL.scala 102:19]
  wire  m_452_io_x2; // @[MUL.scala 102:19]
  wire  m_452_io_x3; // @[MUL.scala 102:19]
  wire  m_452_io_s; // @[MUL.scala 102:19]
  wire  m_452_io_cout; // @[MUL.scala 102:19]
  wire  m_453_io_x1; // @[MUL.scala 102:19]
  wire  m_453_io_x2; // @[MUL.scala 102:19]
  wire  m_453_io_x3; // @[MUL.scala 102:19]
  wire  m_453_io_s; // @[MUL.scala 102:19]
  wire  m_453_io_cout; // @[MUL.scala 102:19]
  wire  m_454_io_x1; // @[MUL.scala 102:19]
  wire  m_454_io_x2; // @[MUL.scala 102:19]
  wire  m_454_io_x3; // @[MUL.scala 102:19]
  wire  m_454_io_s; // @[MUL.scala 102:19]
  wire  m_454_io_cout; // @[MUL.scala 102:19]
  wire  m_455_io_x1; // @[MUL.scala 102:19]
  wire  m_455_io_x2; // @[MUL.scala 102:19]
  wire  m_455_io_x3; // @[MUL.scala 102:19]
  wire  m_455_io_s; // @[MUL.scala 102:19]
  wire  m_455_io_cout; // @[MUL.scala 102:19]
  wire  m_456_io_x1; // @[MUL.scala 102:19]
  wire  m_456_io_x2; // @[MUL.scala 102:19]
  wire  m_456_io_x3; // @[MUL.scala 102:19]
  wire  m_456_io_s; // @[MUL.scala 102:19]
  wire  m_456_io_cout; // @[MUL.scala 102:19]
  wire  m_457_io_x1; // @[MUL.scala 102:19]
  wire  m_457_io_x2; // @[MUL.scala 102:19]
  wire  m_457_io_x3; // @[MUL.scala 102:19]
  wire  m_457_io_s; // @[MUL.scala 102:19]
  wire  m_457_io_cout; // @[MUL.scala 102:19]
  wire  m_458_io_x1; // @[MUL.scala 102:19]
  wire  m_458_io_x2; // @[MUL.scala 102:19]
  wire  m_458_io_x3; // @[MUL.scala 102:19]
  wire  m_458_io_s; // @[MUL.scala 102:19]
  wire  m_458_io_cout; // @[MUL.scala 102:19]
  wire  m_459_io_x1; // @[MUL.scala 102:19]
  wire  m_459_io_x2; // @[MUL.scala 102:19]
  wire  m_459_io_x3; // @[MUL.scala 102:19]
  wire  m_459_io_s; // @[MUL.scala 102:19]
  wire  m_459_io_cout; // @[MUL.scala 102:19]
  wire  m_460_io_x1; // @[MUL.scala 102:19]
  wire  m_460_io_x2; // @[MUL.scala 102:19]
  wire  m_460_io_x3; // @[MUL.scala 102:19]
  wire  m_460_io_s; // @[MUL.scala 102:19]
  wire  m_460_io_cout; // @[MUL.scala 102:19]
  wire  m_461_io_x1; // @[MUL.scala 102:19]
  wire  m_461_io_x2; // @[MUL.scala 102:19]
  wire  m_461_io_x3; // @[MUL.scala 102:19]
  wire  m_461_io_s; // @[MUL.scala 102:19]
  wire  m_461_io_cout; // @[MUL.scala 102:19]
  wire  m_462_io_x1; // @[MUL.scala 102:19]
  wire  m_462_io_x2; // @[MUL.scala 102:19]
  wire  m_462_io_x3; // @[MUL.scala 102:19]
  wire  m_462_io_s; // @[MUL.scala 102:19]
  wire  m_462_io_cout; // @[MUL.scala 102:19]
  wire  m_463_io_x1; // @[MUL.scala 102:19]
  wire  m_463_io_x2; // @[MUL.scala 102:19]
  wire  m_463_io_x3; // @[MUL.scala 102:19]
  wire  m_463_io_s; // @[MUL.scala 102:19]
  wire  m_463_io_cout; // @[MUL.scala 102:19]
  wire  m_464_io_x1; // @[MUL.scala 102:19]
  wire  m_464_io_x2; // @[MUL.scala 102:19]
  wire  m_464_io_x3; // @[MUL.scala 102:19]
  wire  m_464_io_s; // @[MUL.scala 102:19]
  wire  m_464_io_cout; // @[MUL.scala 102:19]
  wire  m_465_io_x1; // @[MUL.scala 102:19]
  wire  m_465_io_x2; // @[MUL.scala 102:19]
  wire  m_465_io_x3; // @[MUL.scala 102:19]
  wire  m_465_io_s; // @[MUL.scala 102:19]
  wire  m_465_io_cout; // @[MUL.scala 102:19]
  wire  m_466_io_x1; // @[MUL.scala 102:19]
  wire  m_466_io_x2; // @[MUL.scala 102:19]
  wire  m_466_io_x3; // @[MUL.scala 102:19]
  wire  m_466_io_s; // @[MUL.scala 102:19]
  wire  m_466_io_cout; // @[MUL.scala 102:19]
  wire  m_467_io_x1; // @[MUL.scala 102:19]
  wire  m_467_io_x2; // @[MUL.scala 102:19]
  wire  m_467_io_x3; // @[MUL.scala 102:19]
  wire  m_467_io_s; // @[MUL.scala 102:19]
  wire  m_467_io_cout; // @[MUL.scala 102:19]
  wire  m_468_io_x1; // @[MUL.scala 102:19]
  wire  m_468_io_x2; // @[MUL.scala 102:19]
  wire  m_468_io_x3; // @[MUL.scala 102:19]
  wire  m_468_io_s; // @[MUL.scala 102:19]
  wire  m_468_io_cout; // @[MUL.scala 102:19]
  wire  m_469_io_x1; // @[MUL.scala 102:19]
  wire  m_469_io_x2; // @[MUL.scala 102:19]
  wire  m_469_io_x3; // @[MUL.scala 102:19]
  wire  m_469_io_s; // @[MUL.scala 102:19]
  wire  m_469_io_cout; // @[MUL.scala 102:19]
  wire  m_470_io_x1; // @[MUL.scala 102:19]
  wire  m_470_io_x2; // @[MUL.scala 102:19]
  wire  m_470_io_x3; // @[MUL.scala 102:19]
  wire  m_470_io_s; // @[MUL.scala 102:19]
  wire  m_470_io_cout; // @[MUL.scala 102:19]
  wire  m_471_io_x1; // @[MUL.scala 102:19]
  wire  m_471_io_x2; // @[MUL.scala 102:19]
  wire  m_471_io_x3; // @[MUL.scala 102:19]
  wire  m_471_io_s; // @[MUL.scala 102:19]
  wire  m_471_io_cout; // @[MUL.scala 102:19]
  wire  m_472_io_in_0; // @[MUL.scala 124:19]
  wire  m_472_io_in_1; // @[MUL.scala 124:19]
  wire  m_472_io_out_0; // @[MUL.scala 124:19]
  wire  m_472_io_out_1; // @[MUL.scala 124:19]
  wire  m_473_io_x1; // @[MUL.scala 102:19]
  wire  m_473_io_x2; // @[MUL.scala 102:19]
  wire  m_473_io_x3; // @[MUL.scala 102:19]
  wire  m_473_io_s; // @[MUL.scala 102:19]
  wire  m_473_io_cout; // @[MUL.scala 102:19]
  wire  m_474_io_x1; // @[MUL.scala 102:19]
  wire  m_474_io_x2; // @[MUL.scala 102:19]
  wire  m_474_io_x3; // @[MUL.scala 102:19]
  wire  m_474_io_s; // @[MUL.scala 102:19]
  wire  m_474_io_cout; // @[MUL.scala 102:19]
  wire  m_475_io_x1; // @[MUL.scala 102:19]
  wire  m_475_io_x2; // @[MUL.scala 102:19]
  wire  m_475_io_x3; // @[MUL.scala 102:19]
  wire  m_475_io_s; // @[MUL.scala 102:19]
  wire  m_475_io_cout; // @[MUL.scala 102:19]
  wire  m_476_io_x1; // @[MUL.scala 102:19]
  wire  m_476_io_x2; // @[MUL.scala 102:19]
  wire  m_476_io_x3; // @[MUL.scala 102:19]
  wire  m_476_io_s; // @[MUL.scala 102:19]
  wire  m_476_io_cout; // @[MUL.scala 102:19]
  wire  m_477_io_x1; // @[MUL.scala 102:19]
  wire  m_477_io_x2; // @[MUL.scala 102:19]
  wire  m_477_io_x3; // @[MUL.scala 102:19]
  wire  m_477_io_s; // @[MUL.scala 102:19]
  wire  m_477_io_cout; // @[MUL.scala 102:19]
  wire  m_478_io_x1; // @[MUL.scala 102:19]
  wire  m_478_io_x2; // @[MUL.scala 102:19]
  wire  m_478_io_x3; // @[MUL.scala 102:19]
  wire  m_478_io_s; // @[MUL.scala 102:19]
  wire  m_478_io_cout; // @[MUL.scala 102:19]
  wire  m_479_io_x1; // @[MUL.scala 102:19]
  wire  m_479_io_x2; // @[MUL.scala 102:19]
  wire  m_479_io_x3; // @[MUL.scala 102:19]
  wire  m_479_io_s; // @[MUL.scala 102:19]
  wire  m_479_io_cout; // @[MUL.scala 102:19]
  wire  m_480_io_x1; // @[MUL.scala 102:19]
  wire  m_480_io_x2; // @[MUL.scala 102:19]
  wire  m_480_io_x3; // @[MUL.scala 102:19]
  wire  m_480_io_s; // @[MUL.scala 102:19]
  wire  m_480_io_cout; // @[MUL.scala 102:19]
  wire  m_481_io_x1; // @[MUL.scala 102:19]
  wire  m_481_io_x2; // @[MUL.scala 102:19]
  wire  m_481_io_x3; // @[MUL.scala 102:19]
  wire  m_481_io_s; // @[MUL.scala 102:19]
  wire  m_481_io_cout; // @[MUL.scala 102:19]
  wire  m_482_io_x1; // @[MUL.scala 102:19]
  wire  m_482_io_x2; // @[MUL.scala 102:19]
  wire  m_482_io_x3; // @[MUL.scala 102:19]
  wire  m_482_io_s; // @[MUL.scala 102:19]
  wire  m_482_io_cout; // @[MUL.scala 102:19]
  wire  m_483_io_x1; // @[MUL.scala 102:19]
  wire  m_483_io_x2; // @[MUL.scala 102:19]
  wire  m_483_io_x3; // @[MUL.scala 102:19]
  wire  m_483_io_s; // @[MUL.scala 102:19]
  wire  m_483_io_cout; // @[MUL.scala 102:19]
  wire  m_484_io_x1; // @[MUL.scala 102:19]
  wire  m_484_io_x2; // @[MUL.scala 102:19]
  wire  m_484_io_x3; // @[MUL.scala 102:19]
  wire  m_484_io_s; // @[MUL.scala 102:19]
  wire  m_484_io_cout; // @[MUL.scala 102:19]
  wire  m_485_io_x1; // @[MUL.scala 102:19]
  wire  m_485_io_x2; // @[MUL.scala 102:19]
  wire  m_485_io_x3; // @[MUL.scala 102:19]
  wire  m_485_io_s; // @[MUL.scala 102:19]
  wire  m_485_io_cout; // @[MUL.scala 102:19]
  wire  m_486_io_x1; // @[MUL.scala 102:19]
  wire  m_486_io_x2; // @[MUL.scala 102:19]
  wire  m_486_io_x3; // @[MUL.scala 102:19]
  wire  m_486_io_s; // @[MUL.scala 102:19]
  wire  m_486_io_cout; // @[MUL.scala 102:19]
  wire  m_487_io_x1; // @[MUL.scala 102:19]
  wire  m_487_io_x2; // @[MUL.scala 102:19]
  wire  m_487_io_x3; // @[MUL.scala 102:19]
  wire  m_487_io_s; // @[MUL.scala 102:19]
  wire  m_487_io_cout; // @[MUL.scala 102:19]
  wire  m_488_io_x1; // @[MUL.scala 102:19]
  wire  m_488_io_x2; // @[MUL.scala 102:19]
  wire  m_488_io_x3; // @[MUL.scala 102:19]
  wire  m_488_io_s; // @[MUL.scala 102:19]
  wire  m_488_io_cout; // @[MUL.scala 102:19]
  wire  m_489_io_x1; // @[MUL.scala 102:19]
  wire  m_489_io_x2; // @[MUL.scala 102:19]
  wire  m_489_io_x3; // @[MUL.scala 102:19]
  wire  m_489_io_s; // @[MUL.scala 102:19]
  wire  m_489_io_cout; // @[MUL.scala 102:19]
  wire  m_490_io_x1; // @[MUL.scala 102:19]
  wire  m_490_io_x2; // @[MUL.scala 102:19]
  wire  m_490_io_x3; // @[MUL.scala 102:19]
  wire  m_490_io_s; // @[MUL.scala 102:19]
  wire  m_490_io_cout; // @[MUL.scala 102:19]
  wire  m_491_io_x1; // @[MUL.scala 102:19]
  wire  m_491_io_x2; // @[MUL.scala 102:19]
  wire  m_491_io_x3; // @[MUL.scala 102:19]
  wire  m_491_io_s; // @[MUL.scala 102:19]
  wire  m_491_io_cout; // @[MUL.scala 102:19]
  wire  m_492_io_x1; // @[MUL.scala 102:19]
  wire  m_492_io_x2; // @[MUL.scala 102:19]
  wire  m_492_io_x3; // @[MUL.scala 102:19]
  wire  m_492_io_s; // @[MUL.scala 102:19]
  wire  m_492_io_cout; // @[MUL.scala 102:19]
  wire  m_493_io_x1; // @[MUL.scala 102:19]
  wire  m_493_io_x2; // @[MUL.scala 102:19]
  wire  m_493_io_x3; // @[MUL.scala 102:19]
  wire  m_493_io_s; // @[MUL.scala 102:19]
  wire  m_493_io_cout; // @[MUL.scala 102:19]
  wire  m_494_io_x1; // @[MUL.scala 102:19]
  wire  m_494_io_x2; // @[MUL.scala 102:19]
  wire  m_494_io_x3; // @[MUL.scala 102:19]
  wire  m_494_io_s; // @[MUL.scala 102:19]
  wire  m_494_io_cout; // @[MUL.scala 102:19]
  wire  m_495_io_x1; // @[MUL.scala 102:19]
  wire  m_495_io_x2; // @[MUL.scala 102:19]
  wire  m_495_io_x3; // @[MUL.scala 102:19]
  wire  m_495_io_s; // @[MUL.scala 102:19]
  wire  m_495_io_cout; // @[MUL.scala 102:19]
  wire  m_496_io_x1; // @[MUL.scala 102:19]
  wire  m_496_io_x2; // @[MUL.scala 102:19]
  wire  m_496_io_x3; // @[MUL.scala 102:19]
  wire  m_496_io_s; // @[MUL.scala 102:19]
  wire  m_496_io_cout; // @[MUL.scala 102:19]
  wire  m_497_io_x1; // @[MUL.scala 102:19]
  wire  m_497_io_x2; // @[MUL.scala 102:19]
  wire  m_497_io_x3; // @[MUL.scala 102:19]
  wire  m_497_io_s; // @[MUL.scala 102:19]
  wire  m_497_io_cout; // @[MUL.scala 102:19]
  wire  m_498_io_x1; // @[MUL.scala 102:19]
  wire  m_498_io_x2; // @[MUL.scala 102:19]
  wire  m_498_io_x3; // @[MUL.scala 102:19]
  wire  m_498_io_s; // @[MUL.scala 102:19]
  wire  m_498_io_cout; // @[MUL.scala 102:19]
  wire  m_499_io_x1; // @[MUL.scala 102:19]
  wire  m_499_io_x2; // @[MUL.scala 102:19]
  wire  m_499_io_x3; // @[MUL.scala 102:19]
  wire  m_499_io_s; // @[MUL.scala 102:19]
  wire  m_499_io_cout; // @[MUL.scala 102:19]
  wire  m_500_io_x1; // @[MUL.scala 102:19]
  wire  m_500_io_x2; // @[MUL.scala 102:19]
  wire  m_500_io_x3; // @[MUL.scala 102:19]
  wire  m_500_io_s; // @[MUL.scala 102:19]
  wire  m_500_io_cout; // @[MUL.scala 102:19]
  wire  m_501_io_x1; // @[MUL.scala 102:19]
  wire  m_501_io_x2; // @[MUL.scala 102:19]
  wire  m_501_io_x3; // @[MUL.scala 102:19]
  wire  m_501_io_s; // @[MUL.scala 102:19]
  wire  m_501_io_cout; // @[MUL.scala 102:19]
  wire  m_502_io_x1; // @[MUL.scala 102:19]
  wire  m_502_io_x2; // @[MUL.scala 102:19]
  wire  m_502_io_x3; // @[MUL.scala 102:19]
  wire  m_502_io_s; // @[MUL.scala 102:19]
  wire  m_502_io_cout; // @[MUL.scala 102:19]
  wire  m_503_io_x1; // @[MUL.scala 102:19]
  wire  m_503_io_x2; // @[MUL.scala 102:19]
  wire  m_503_io_x3; // @[MUL.scala 102:19]
  wire  m_503_io_s; // @[MUL.scala 102:19]
  wire  m_503_io_cout; // @[MUL.scala 102:19]
  wire  m_504_io_x1; // @[MUL.scala 102:19]
  wire  m_504_io_x2; // @[MUL.scala 102:19]
  wire  m_504_io_x3; // @[MUL.scala 102:19]
  wire  m_504_io_s; // @[MUL.scala 102:19]
  wire  m_504_io_cout; // @[MUL.scala 102:19]
  wire  m_505_io_x1; // @[MUL.scala 102:19]
  wire  m_505_io_x2; // @[MUL.scala 102:19]
  wire  m_505_io_x3; // @[MUL.scala 102:19]
  wire  m_505_io_s; // @[MUL.scala 102:19]
  wire  m_505_io_cout; // @[MUL.scala 102:19]
  wire  m_506_io_x1; // @[MUL.scala 102:19]
  wire  m_506_io_x2; // @[MUL.scala 102:19]
  wire  m_506_io_x3; // @[MUL.scala 102:19]
  wire  m_506_io_s; // @[MUL.scala 102:19]
  wire  m_506_io_cout; // @[MUL.scala 102:19]
  wire  m_507_io_x1; // @[MUL.scala 102:19]
  wire  m_507_io_x2; // @[MUL.scala 102:19]
  wire  m_507_io_x3; // @[MUL.scala 102:19]
  wire  m_507_io_s; // @[MUL.scala 102:19]
  wire  m_507_io_cout; // @[MUL.scala 102:19]
  wire  m_508_io_x1; // @[MUL.scala 102:19]
  wire  m_508_io_x2; // @[MUL.scala 102:19]
  wire  m_508_io_x3; // @[MUL.scala 102:19]
  wire  m_508_io_s; // @[MUL.scala 102:19]
  wire  m_508_io_cout; // @[MUL.scala 102:19]
  wire  m_509_io_x1; // @[MUL.scala 102:19]
  wire  m_509_io_x2; // @[MUL.scala 102:19]
  wire  m_509_io_x3; // @[MUL.scala 102:19]
  wire  m_509_io_s; // @[MUL.scala 102:19]
  wire  m_509_io_cout; // @[MUL.scala 102:19]
  wire  m_510_io_x1; // @[MUL.scala 102:19]
  wire  m_510_io_x2; // @[MUL.scala 102:19]
  wire  m_510_io_x3; // @[MUL.scala 102:19]
  wire  m_510_io_s; // @[MUL.scala 102:19]
  wire  m_510_io_cout; // @[MUL.scala 102:19]
  wire  m_511_io_x1; // @[MUL.scala 102:19]
  wire  m_511_io_x2; // @[MUL.scala 102:19]
  wire  m_511_io_x3; // @[MUL.scala 102:19]
  wire  m_511_io_s; // @[MUL.scala 102:19]
  wire  m_511_io_cout; // @[MUL.scala 102:19]
  wire  m_512_io_x1; // @[MUL.scala 102:19]
  wire  m_512_io_x2; // @[MUL.scala 102:19]
  wire  m_512_io_x3; // @[MUL.scala 102:19]
  wire  m_512_io_s; // @[MUL.scala 102:19]
  wire  m_512_io_cout; // @[MUL.scala 102:19]
  wire  m_513_io_x1; // @[MUL.scala 102:19]
  wire  m_513_io_x2; // @[MUL.scala 102:19]
  wire  m_513_io_x3; // @[MUL.scala 102:19]
  wire  m_513_io_s; // @[MUL.scala 102:19]
  wire  m_513_io_cout; // @[MUL.scala 102:19]
  wire  m_514_io_x1; // @[MUL.scala 102:19]
  wire  m_514_io_x2; // @[MUL.scala 102:19]
  wire  m_514_io_x3; // @[MUL.scala 102:19]
  wire  m_514_io_s; // @[MUL.scala 102:19]
  wire  m_514_io_cout; // @[MUL.scala 102:19]
  wire  m_515_io_x1; // @[MUL.scala 102:19]
  wire  m_515_io_x2; // @[MUL.scala 102:19]
  wire  m_515_io_x3; // @[MUL.scala 102:19]
  wire  m_515_io_s; // @[MUL.scala 102:19]
  wire  m_515_io_cout; // @[MUL.scala 102:19]
  wire  m_516_io_x1; // @[MUL.scala 102:19]
  wire  m_516_io_x2; // @[MUL.scala 102:19]
  wire  m_516_io_x3; // @[MUL.scala 102:19]
  wire  m_516_io_s; // @[MUL.scala 102:19]
  wire  m_516_io_cout; // @[MUL.scala 102:19]
  wire  m_517_io_x1; // @[MUL.scala 102:19]
  wire  m_517_io_x2; // @[MUL.scala 102:19]
  wire  m_517_io_x3; // @[MUL.scala 102:19]
  wire  m_517_io_s; // @[MUL.scala 102:19]
  wire  m_517_io_cout; // @[MUL.scala 102:19]
  wire  m_518_io_x1; // @[MUL.scala 102:19]
  wire  m_518_io_x2; // @[MUL.scala 102:19]
  wire  m_518_io_x3; // @[MUL.scala 102:19]
  wire  m_518_io_s; // @[MUL.scala 102:19]
  wire  m_518_io_cout; // @[MUL.scala 102:19]
  wire  m_519_io_x1; // @[MUL.scala 102:19]
  wire  m_519_io_x2; // @[MUL.scala 102:19]
  wire  m_519_io_x3; // @[MUL.scala 102:19]
  wire  m_519_io_s; // @[MUL.scala 102:19]
  wire  m_519_io_cout; // @[MUL.scala 102:19]
  wire  m_520_io_x1; // @[MUL.scala 102:19]
  wire  m_520_io_x2; // @[MUL.scala 102:19]
  wire  m_520_io_x3; // @[MUL.scala 102:19]
  wire  m_520_io_s; // @[MUL.scala 102:19]
  wire  m_520_io_cout; // @[MUL.scala 102:19]
  wire  m_521_io_x1; // @[MUL.scala 102:19]
  wire  m_521_io_x2; // @[MUL.scala 102:19]
  wire  m_521_io_x3; // @[MUL.scala 102:19]
  wire  m_521_io_s; // @[MUL.scala 102:19]
  wire  m_521_io_cout; // @[MUL.scala 102:19]
  wire  m_522_io_in_0; // @[MUL.scala 124:19]
  wire  m_522_io_in_1; // @[MUL.scala 124:19]
  wire  m_522_io_out_0; // @[MUL.scala 124:19]
  wire  m_522_io_out_1; // @[MUL.scala 124:19]
  wire  m_523_io_x1; // @[MUL.scala 102:19]
  wire  m_523_io_x2; // @[MUL.scala 102:19]
  wire  m_523_io_x3; // @[MUL.scala 102:19]
  wire  m_523_io_s; // @[MUL.scala 102:19]
  wire  m_523_io_cout; // @[MUL.scala 102:19]
  wire  m_524_io_x1; // @[MUL.scala 102:19]
  wire  m_524_io_x2; // @[MUL.scala 102:19]
  wire  m_524_io_x3; // @[MUL.scala 102:19]
  wire  m_524_io_s; // @[MUL.scala 102:19]
  wire  m_524_io_cout; // @[MUL.scala 102:19]
  wire  m_525_io_x1; // @[MUL.scala 102:19]
  wire  m_525_io_x2; // @[MUL.scala 102:19]
  wire  m_525_io_x3; // @[MUL.scala 102:19]
  wire  m_525_io_s; // @[MUL.scala 102:19]
  wire  m_525_io_cout; // @[MUL.scala 102:19]
  wire  m_526_io_x1; // @[MUL.scala 102:19]
  wire  m_526_io_x2; // @[MUL.scala 102:19]
  wire  m_526_io_x3; // @[MUL.scala 102:19]
  wire  m_526_io_s; // @[MUL.scala 102:19]
  wire  m_526_io_cout; // @[MUL.scala 102:19]
  wire  m_527_io_x1; // @[MUL.scala 102:19]
  wire  m_527_io_x2; // @[MUL.scala 102:19]
  wire  m_527_io_x3; // @[MUL.scala 102:19]
  wire  m_527_io_s; // @[MUL.scala 102:19]
  wire  m_527_io_cout; // @[MUL.scala 102:19]
  wire  m_528_io_x1; // @[MUL.scala 102:19]
  wire  m_528_io_x2; // @[MUL.scala 102:19]
  wire  m_528_io_x3; // @[MUL.scala 102:19]
  wire  m_528_io_s; // @[MUL.scala 102:19]
  wire  m_528_io_cout; // @[MUL.scala 102:19]
  wire  m_529_io_x1; // @[MUL.scala 102:19]
  wire  m_529_io_x2; // @[MUL.scala 102:19]
  wire  m_529_io_x3; // @[MUL.scala 102:19]
  wire  m_529_io_s; // @[MUL.scala 102:19]
  wire  m_529_io_cout; // @[MUL.scala 102:19]
  wire  m_530_io_x1; // @[MUL.scala 102:19]
  wire  m_530_io_x2; // @[MUL.scala 102:19]
  wire  m_530_io_x3; // @[MUL.scala 102:19]
  wire  m_530_io_s; // @[MUL.scala 102:19]
  wire  m_530_io_cout; // @[MUL.scala 102:19]
  wire  m_531_io_x1; // @[MUL.scala 102:19]
  wire  m_531_io_x2; // @[MUL.scala 102:19]
  wire  m_531_io_x3; // @[MUL.scala 102:19]
  wire  m_531_io_s; // @[MUL.scala 102:19]
  wire  m_531_io_cout; // @[MUL.scala 102:19]
  wire  m_532_io_in_0; // @[MUL.scala 124:19]
  wire  m_532_io_in_1; // @[MUL.scala 124:19]
  wire  m_532_io_out_0; // @[MUL.scala 124:19]
  wire  m_532_io_out_1; // @[MUL.scala 124:19]
  wire  m_533_io_x1; // @[MUL.scala 102:19]
  wire  m_533_io_x2; // @[MUL.scala 102:19]
  wire  m_533_io_x3; // @[MUL.scala 102:19]
  wire  m_533_io_s; // @[MUL.scala 102:19]
  wire  m_533_io_cout; // @[MUL.scala 102:19]
  wire  m_534_io_x1; // @[MUL.scala 102:19]
  wire  m_534_io_x2; // @[MUL.scala 102:19]
  wire  m_534_io_x3; // @[MUL.scala 102:19]
  wire  m_534_io_s; // @[MUL.scala 102:19]
  wire  m_534_io_cout; // @[MUL.scala 102:19]
  wire  m_535_io_x1; // @[MUL.scala 102:19]
  wire  m_535_io_x2; // @[MUL.scala 102:19]
  wire  m_535_io_x3; // @[MUL.scala 102:19]
  wire  m_535_io_s; // @[MUL.scala 102:19]
  wire  m_535_io_cout; // @[MUL.scala 102:19]
  wire  m_536_io_x1; // @[MUL.scala 102:19]
  wire  m_536_io_x2; // @[MUL.scala 102:19]
  wire  m_536_io_x3; // @[MUL.scala 102:19]
  wire  m_536_io_s; // @[MUL.scala 102:19]
  wire  m_536_io_cout; // @[MUL.scala 102:19]
  wire  m_537_io_x1; // @[MUL.scala 102:19]
  wire  m_537_io_x2; // @[MUL.scala 102:19]
  wire  m_537_io_x3; // @[MUL.scala 102:19]
  wire  m_537_io_s; // @[MUL.scala 102:19]
  wire  m_537_io_cout; // @[MUL.scala 102:19]
  wire  m_538_io_x1; // @[MUL.scala 102:19]
  wire  m_538_io_x2; // @[MUL.scala 102:19]
  wire  m_538_io_x3; // @[MUL.scala 102:19]
  wire  m_538_io_s; // @[MUL.scala 102:19]
  wire  m_538_io_cout; // @[MUL.scala 102:19]
  wire  m_539_io_x1; // @[MUL.scala 102:19]
  wire  m_539_io_x2; // @[MUL.scala 102:19]
  wire  m_539_io_x3; // @[MUL.scala 102:19]
  wire  m_539_io_s; // @[MUL.scala 102:19]
  wire  m_539_io_cout; // @[MUL.scala 102:19]
  wire  m_540_io_x1; // @[MUL.scala 102:19]
  wire  m_540_io_x2; // @[MUL.scala 102:19]
  wire  m_540_io_x3; // @[MUL.scala 102:19]
  wire  m_540_io_s; // @[MUL.scala 102:19]
  wire  m_540_io_cout; // @[MUL.scala 102:19]
  wire  m_541_io_x1; // @[MUL.scala 102:19]
  wire  m_541_io_x2; // @[MUL.scala 102:19]
  wire  m_541_io_x3; // @[MUL.scala 102:19]
  wire  m_541_io_s; // @[MUL.scala 102:19]
  wire  m_541_io_cout; // @[MUL.scala 102:19]
  wire  m_542_io_x1; // @[MUL.scala 102:19]
  wire  m_542_io_x2; // @[MUL.scala 102:19]
  wire  m_542_io_x3; // @[MUL.scala 102:19]
  wire  m_542_io_s; // @[MUL.scala 102:19]
  wire  m_542_io_cout; // @[MUL.scala 102:19]
  wire  m_543_io_x1; // @[MUL.scala 102:19]
  wire  m_543_io_x2; // @[MUL.scala 102:19]
  wire  m_543_io_x3; // @[MUL.scala 102:19]
  wire  m_543_io_s; // @[MUL.scala 102:19]
  wire  m_543_io_cout; // @[MUL.scala 102:19]
  wire  m_544_io_x1; // @[MUL.scala 102:19]
  wire  m_544_io_x2; // @[MUL.scala 102:19]
  wire  m_544_io_x3; // @[MUL.scala 102:19]
  wire  m_544_io_s; // @[MUL.scala 102:19]
  wire  m_544_io_cout; // @[MUL.scala 102:19]
  wire  m_545_io_x1; // @[MUL.scala 102:19]
  wire  m_545_io_x2; // @[MUL.scala 102:19]
  wire  m_545_io_x3; // @[MUL.scala 102:19]
  wire  m_545_io_s; // @[MUL.scala 102:19]
  wire  m_545_io_cout; // @[MUL.scala 102:19]
  wire  m_546_io_x1; // @[MUL.scala 102:19]
  wire  m_546_io_x2; // @[MUL.scala 102:19]
  wire  m_546_io_x3; // @[MUL.scala 102:19]
  wire  m_546_io_s; // @[MUL.scala 102:19]
  wire  m_546_io_cout; // @[MUL.scala 102:19]
  wire  m_547_io_x1; // @[MUL.scala 102:19]
  wire  m_547_io_x2; // @[MUL.scala 102:19]
  wire  m_547_io_x3; // @[MUL.scala 102:19]
  wire  m_547_io_s; // @[MUL.scala 102:19]
  wire  m_547_io_cout; // @[MUL.scala 102:19]
  wire  m_548_io_x1; // @[MUL.scala 102:19]
  wire  m_548_io_x2; // @[MUL.scala 102:19]
  wire  m_548_io_x3; // @[MUL.scala 102:19]
  wire  m_548_io_s; // @[MUL.scala 102:19]
  wire  m_548_io_cout; // @[MUL.scala 102:19]
  wire  m_549_io_x1; // @[MUL.scala 102:19]
  wire  m_549_io_x2; // @[MUL.scala 102:19]
  wire  m_549_io_x3; // @[MUL.scala 102:19]
  wire  m_549_io_s; // @[MUL.scala 102:19]
  wire  m_549_io_cout; // @[MUL.scala 102:19]
  wire  m_550_io_x1; // @[MUL.scala 102:19]
  wire  m_550_io_x2; // @[MUL.scala 102:19]
  wire  m_550_io_x3; // @[MUL.scala 102:19]
  wire  m_550_io_s; // @[MUL.scala 102:19]
  wire  m_550_io_cout; // @[MUL.scala 102:19]
  wire  m_551_io_x1; // @[MUL.scala 102:19]
  wire  m_551_io_x2; // @[MUL.scala 102:19]
  wire  m_551_io_x3; // @[MUL.scala 102:19]
  wire  m_551_io_s; // @[MUL.scala 102:19]
  wire  m_551_io_cout; // @[MUL.scala 102:19]
  wire  m_552_io_x1; // @[MUL.scala 102:19]
  wire  m_552_io_x2; // @[MUL.scala 102:19]
  wire  m_552_io_x3; // @[MUL.scala 102:19]
  wire  m_552_io_s; // @[MUL.scala 102:19]
  wire  m_552_io_cout; // @[MUL.scala 102:19]
  wire  m_553_io_x1; // @[MUL.scala 102:19]
  wire  m_553_io_x2; // @[MUL.scala 102:19]
  wire  m_553_io_x3; // @[MUL.scala 102:19]
  wire  m_553_io_s; // @[MUL.scala 102:19]
  wire  m_553_io_cout; // @[MUL.scala 102:19]
  wire  m_554_io_x1; // @[MUL.scala 102:19]
  wire  m_554_io_x2; // @[MUL.scala 102:19]
  wire  m_554_io_x3; // @[MUL.scala 102:19]
  wire  m_554_io_s; // @[MUL.scala 102:19]
  wire  m_554_io_cout; // @[MUL.scala 102:19]
  wire  m_555_io_x1; // @[MUL.scala 102:19]
  wire  m_555_io_x2; // @[MUL.scala 102:19]
  wire  m_555_io_x3; // @[MUL.scala 102:19]
  wire  m_555_io_s; // @[MUL.scala 102:19]
  wire  m_555_io_cout; // @[MUL.scala 102:19]
  wire  m_556_io_x1; // @[MUL.scala 102:19]
  wire  m_556_io_x2; // @[MUL.scala 102:19]
  wire  m_556_io_x3; // @[MUL.scala 102:19]
  wire  m_556_io_s; // @[MUL.scala 102:19]
  wire  m_556_io_cout; // @[MUL.scala 102:19]
  wire  m_557_io_x1; // @[MUL.scala 102:19]
  wire  m_557_io_x2; // @[MUL.scala 102:19]
  wire  m_557_io_x3; // @[MUL.scala 102:19]
  wire  m_557_io_s; // @[MUL.scala 102:19]
  wire  m_557_io_cout; // @[MUL.scala 102:19]
  wire  m_558_io_x1; // @[MUL.scala 102:19]
  wire  m_558_io_x2; // @[MUL.scala 102:19]
  wire  m_558_io_x3; // @[MUL.scala 102:19]
  wire  m_558_io_s; // @[MUL.scala 102:19]
  wire  m_558_io_cout; // @[MUL.scala 102:19]
  wire  m_559_io_x1; // @[MUL.scala 102:19]
  wire  m_559_io_x2; // @[MUL.scala 102:19]
  wire  m_559_io_x3; // @[MUL.scala 102:19]
  wire  m_559_io_s; // @[MUL.scala 102:19]
  wire  m_559_io_cout; // @[MUL.scala 102:19]
  wire  m_560_io_x1; // @[MUL.scala 102:19]
  wire  m_560_io_x2; // @[MUL.scala 102:19]
  wire  m_560_io_x3; // @[MUL.scala 102:19]
  wire  m_560_io_s; // @[MUL.scala 102:19]
  wire  m_560_io_cout; // @[MUL.scala 102:19]
  wire  m_561_io_x1; // @[MUL.scala 102:19]
  wire  m_561_io_x2; // @[MUL.scala 102:19]
  wire  m_561_io_x3; // @[MUL.scala 102:19]
  wire  m_561_io_s; // @[MUL.scala 102:19]
  wire  m_561_io_cout; // @[MUL.scala 102:19]
  wire  m_562_io_x1; // @[MUL.scala 102:19]
  wire  m_562_io_x2; // @[MUL.scala 102:19]
  wire  m_562_io_x3; // @[MUL.scala 102:19]
  wire  m_562_io_s; // @[MUL.scala 102:19]
  wire  m_562_io_cout; // @[MUL.scala 102:19]
  wire  m_563_io_x1; // @[MUL.scala 102:19]
  wire  m_563_io_x2; // @[MUL.scala 102:19]
  wire  m_563_io_x3; // @[MUL.scala 102:19]
  wire  m_563_io_s; // @[MUL.scala 102:19]
  wire  m_563_io_cout; // @[MUL.scala 102:19]
  wire  m_564_io_x1; // @[MUL.scala 102:19]
  wire  m_564_io_x2; // @[MUL.scala 102:19]
  wire  m_564_io_x3; // @[MUL.scala 102:19]
  wire  m_564_io_s; // @[MUL.scala 102:19]
  wire  m_564_io_cout; // @[MUL.scala 102:19]
  wire  m_565_io_x1; // @[MUL.scala 102:19]
  wire  m_565_io_x2; // @[MUL.scala 102:19]
  wire  m_565_io_x3; // @[MUL.scala 102:19]
  wire  m_565_io_s; // @[MUL.scala 102:19]
  wire  m_565_io_cout; // @[MUL.scala 102:19]
  wire  m_566_io_x1; // @[MUL.scala 102:19]
  wire  m_566_io_x2; // @[MUL.scala 102:19]
  wire  m_566_io_x3; // @[MUL.scala 102:19]
  wire  m_566_io_s; // @[MUL.scala 102:19]
  wire  m_566_io_cout; // @[MUL.scala 102:19]
  wire  m_567_io_x1; // @[MUL.scala 102:19]
  wire  m_567_io_x2; // @[MUL.scala 102:19]
  wire  m_567_io_x3; // @[MUL.scala 102:19]
  wire  m_567_io_s; // @[MUL.scala 102:19]
  wire  m_567_io_cout; // @[MUL.scala 102:19]
  wire  m_568_io_x1; // @[MUL.scala 102:19]
  wire  m_568_io_x2; // @[MUL.scala 102:19]
  wire  m_568_io_x3; // @[MUL.scala 102:19]
  wire  m_568_io_s; // @[MUL.scala 102:19]
  wire  m_568_io_cout; // @[MUL.scala 102:19]
  wire  m_569_io_x1; // @[MUL.scala 102:19]
  wire  m_569_io_x2; // @[MUL.scala 102:19]
  wire  m_569_io_x3; // @[MUL.scala 102:19]
  wire  m_569_io_s; // @[MUL.scala 102:19]
  wire  m_569_io_cout; // @[MUL.scala 102:19]
  wire  m_570_io_x1; // @[MUL.scala 102:19]
  wire  m_570_io_x2; // @[MUL.scala 102:19]
  wire  m_570_io_x3; // @[MUL.scala 102:19]
  wire  m_570_io_s; // @[MUL.scala 102:19]
  wire  m_570_io_cout; // @[MUL.scala 102:19]
  wire  m_571_io_x1; // @[MUL.scala 102:19]
  wire  m_571_io_x2; // @[MUL.scala 102:19]
  wire  m_571_io_x3; // @[MUL.scala 102:19]
  wire  m_571_io_s; // @[MUL.scala 102:19]
  wire  m_571_io_cout; // @[MUL.scala 102:19]
  wire  m_572_io_x1; // @[MUL.scala 102:19]
  wire  m_572_io_x2; // @[MUL.scala 102:19]
  wire  m_572_io_x3; // @[MUL.scala 102:19]
  wire  m_572_io_s; // @[MUL.scala 102:19]
  wire  m_572_io_cout; // @[MUL.scala 102:19]
  wire  m_573_io_x1; // @[MUL.scala 102:19]
  wire  m_573_io_x2; // @[MUL.scala 102:19]
  wire  m_573_io_x3; // @[MUL.scala 102:19]
  wire  m_573_io_s; // @[MUL.scala 102:19]
  wire  m_573_io_cout; // @[MUL.scala 102:19]
  wire  m_574_io_x1; // @[MUL.scala 102:19]
  wire  m_574_io_x2; // @[MUL.scala 102:19]
  wire  m_574_io_x3; // @[MUL.scala 102:19]
  wire  m_574_io_s; // @[MUL.scala 102:19]
  wire  m_574_io_cout; // @[MUL.scala 102:19]
  wire  m_575_io_x1; // @[MUL.scala 102:19]
  wire  m_575_io_x2; // @[MUL.scala 102:19]
  wire  m_575_io_x3; // @[MUL.scala 102:19]
  wire  m_575_io_s; // @[MUL.scala 102:19]
  wire  m_575_io_cout; // @[MUL.scala 102:19]
  wire  m_576_io_x1; // @[MUL.scala 102:19]
  wire  m_576_io_x2; // @[MUL.scala 102:19]
  wire  m_576_io_x3; // @[MUL.scala 102:19]
  wire  m_576_io_s; // @[MUL.scala 102:19]
  wire  m_576_io_cout; // @[MUL.scala 102:19]
  wire  m_577_io_in_0; // @[MUL.scala 124:19]
  wire  m_577_io_in_1; // @[MUL.scala 124:19]
  wire  m_577_io_out_0; // @[MUL.scala 124:19]
  wire  m_577_io_out_1; // @[MUL.scala 124:19]
  wire  m_578_io_x1; // @[MUL.scala 102:19]
  wire  m_578_io_x2; // @[MUL.scala 102:19]
  wire  m_578_io_x3; // @[MUL.scala 102:19]
  wire  m_578_io_s; // @[MUL.scala 102:19]
  wire  m_578_io_cout; // @[MUL.scala 102:19]
  wire  m_579_io_x1; // @[MUL.scala 102:19]
  wire  m_579_io_x2; // @[MUL.scala 102:19]
  wire  m_579_io_x3; // @[MUL.scala 102:19]
  wire  m_579_io_s; // @[MUL.scala 102:19]
  wire  m_579_io_cout; // @[MUL.scala 102:19]
  wire  m_580_io_x1; // @[MUL.scala 102:19]
  wire  m_580_io_x2; // @[MUL.scala 102:19]
  wire  m_580_io_x3; // @[MUL.scala 102:19]
  wire  m_580_io_s; // @[MUL.scala 102:19]
  wire  m_580_io_cout; // @[MUL.scala 102:19]
  wire  m_581_io_x1; // @[MUL.scala 102:19]
  wire  m_581_io_x2; // @[MUL.scala 102:19]
  wire  m_581_io_x3; // @[MUL.scala 102:19]
  wire  m_581_io_s; // @[MUL.scala 102:19]
  wire  m_581_io_cout; // @[MUL.scala 102:19]
  wire  m_582_io_x1; // @[MUL.scala 102:19]
  wire  m_582_io_x2; // @[MUL.scala 102:19]
  wire  m_582_io_x3; // @[MUL.scala 102:19]
  wire  m_582_io_s; // @[MUL.scala 102:19]
  wire  m_582_io_cout; // @[MUL.scala 102:19]
  wire  m_583_io_x1; // @[MUL.scala 102:19]
  wire  m_583_io_x2; // @[MUL.scala 102:19]
  wire  m_583_io_x3; // @[MUL.scala 102:19]
  wire  m_583_io_s; // @[MUL.scala 102:19]
  wire  m_583_io_cout; // @[MUL.scala 102:19]
  wire  m_584_io_x1; // @[MUL.scala 102:19]
  wire  m_584_io_x2; // @[MUL.scala 102:19]
  wire  m_584_io_x3; // @[MUL.scala 102:19]
  wire  m_584_io_s; // @[MUL.scala 102:19]
  wire  m_584_io_cout; // @[MUL.scala 102:19]
  wire  m_585_io_x1; // @[MUL.scala 102:19]
  wire  m_585_io_x2; // @[MUL.scala 102:19]
  wire  m_585_io_x3; // @[MUL.scala 102:19]
  wire  m_585_io_s; // @[MUL.scala 102:19]
  wire  m_585_io_cout; // @[MUL.scala 102:19]
  wire  m_586_io_in_0; // @[MUL.scala 124:19]
  wire  m_586_io_in_1; // @[MUL.scala 124:19]
  wire  m_586_io_out_0; // @[MUL.scala 124:19]
  wire  m_586_io_out_1; // @[MUL.scala 124:19]
  wire  m_587_io_x1; // @[MUL.scala 102:19]
  wire  m_587_io_x2; // @[MUL.scala 102:19]
  wire  m_587_io_x3; // @[MUL.scala 102:19]
  wire  m_587_io_s; // @[MUL.scala 102:19]
  wire  m_587_io_cout; // @[MUL.scala 102:19]
  wire  m_588_io_x1; // @[MUL.scala 102:19]
  wire  m_588_io_x2; // @[MUL.scala 102:19]
  wire  m_588_io_x3; // @[MUL.scala 102:19]
  wire  m_588_io_s; // @[MUL.scala 102:19]
  wire  m_588_io_cout; // @[MUL.scala 102:19]
  wire  m_589_io_x1; // @[MUL.scala 102:19]
  wire  m_589_io_x2; // @[MUL.scala 102:19]
  wire  m_589_io_x3; // @[MUL.scala 102:19]
  wire  m_589_io_s; // @[MUL.scala 102:19]
  wire  m_589_io_cout; // @[MUL.scala 102:19]
  wire  m_590_io_x1; // @[MUL.scala 102:19]
  wire  m_590_io_x2; // @[MUL.scala 102:19]
  wire  m_590_io_x3; // @[MUL.scala 102:19]
  wire  m_590_io_s; // @[MUL.scala 102:19]
  wire  m_590_io_cout; // @[MUL.scala 102:19]
  wire  m_591_io_x1; // @[MUL.scala 102:19]
  wire  m_591_io_x2; // @[MUL.scala 102:19]
  wire  m_591_io_x3; // @[MUL.scala 102:19]
  wire  m_591_io_s; // @[MUL.scala 102:19]
  wire  m_591_io_cout; // @[MUL.scala 102:19]
  wire  m_592_io_x1; // @[MUL.scala 102:19]
  wire  m_592_io_x2; // @[MUL.scala 102:19]
  wire  m_592_io_x3; // @[MUL.scala 102:19]
  wire  m_592_io_s; // @[MUL.scala 102:19]
  wire  m_592_io_cout; // @[MUL.scala 102:19]
  wire  m_593_io_x1; // @[MUL.scala 102:19]
  wire  m_593_io_x2; // @[MUL.scala 102:19]
  wire  m_593_io_x3; // @[MUL.scala 102:19]
  wire  m_593_io_s; // @[MUL.scala 102:19]
  wire  m_593_io_cout; // @[MUL.scala 102:19]
  wire  m_594_io_x1; // @[MUL.scala 102:19]
  wire  m_594_io_x2; // @[MUL.scala 102:19]
  wire  m_594_io_x3; // @[MUL.scala 102:19]
  wire  m_594_io_s; // @[MUL.scala 102:19]
  wire  m_594_io_cout; // @[MUL.scala 102:19]
  wire  m_595_io_x1; // @[MUL.scala 102:19]
  wire  m_595_io_x2; // @[MUL.scala 102:19]
  wire  m_595_io_x3; // @[MUL.scala 102:19]
  wire  m_595_io_s; // @[MUL.scala 102:19]
  wire  m_595_io_cout; // @[MUL.scala 102:19]
  wire  m_596_io_x1; // @[MUL.scala 102:19]
  wire  m_596_io_x2; // @[MUL.scala 102:19]
  wire  m_596_io_x3; // @[MUL.scala 102:19]
  wire  m_596_io_s; // @[MUL.scala 102:19]
  wire  m_596_io_cout; // @[MUL.scala 102:19]
  wire  m_597_io_x1; // @[MUL.scala 102:19]
  wire  m_597_io_x2; // @[MUL.scala 102:19]
  wire  m_597_io_x3; // @[MUL.scala 102:19]
  wire  m_597_io_s; // @[MUL.scala 102:19]
  wire  m_597_io_cout; // @[MUL.scala 102:19]
  wire  m_598_io_x1; // @[MUL.scala 102:19]
  wire  m_598_io_x2; // @[MUL.scala 102:19]
  wire  m_598_io_x3; // @[MUL.scala 102:19]
  wire  m_598_io_s; // @[MUL.scala 102:19]
  wire  m_598_io_cout; // @[MUL.scala 102:19]
  wire  m_599_io_x1; // @[MUL.scala 102:19]
  wire  m_599_io_x2; // @[MUL.scala 102:19]
  wire  m_599_io_x3; // @[MUL.scala 102:19]
  wire  m_599_io_s; // @[MUL.scala 102:19]
  wire  m_599_io_cout; // @[MUL.scala 102:19]
  wire  m_600_io_x1; // @[MUL.scala 102:19]
  wire  m_600_io_x2; // @[MUL.scala 102:19]
  wire  m_600_io_x3; // @[MUL.scala 102:19]
  wire  m_600_io_s; // @[MUL.scala 102:19]
  wire  m_600_io_cout; // @[MUL.scala 102:19]
  wire  m_601_io_x1; // @[MUL.scala 102:19]
  wire  m_601_io_x2; // @[MUL.scala 102:19]
  wire  m_601_io_x3; // @[MUL.scala 102:19]
  wire  m_601_io_s; // @[MUL.scala 102:19]
  wire  m_601_io_cout; // @[MUL.scala 102:19]
  wire  m_602_io_x1; // @[MUL.scala 102:19]
  wire  m_602_io_x2; // @[MUL.scala 102:19]
  wire  m_602_io_x3; // @[MUL.scala 102:19]
  wire  m_602_io_s; // @[MUL.scala 102:19]
  wire  m_602_io_cout; // @[MUL.scala 102:19]
  wire  m_603_io_x1; // @[MUL.scala 102:19]
  wire  m_603_io_x2; // @[MUL.scala 102:19]
  wire  m_603_io_x3; // @[MUL.scala 102:19]
  wire  m_603_io_s; // @[MUL.scala 102:19]
  wire  m_603_io_cout; // @[MUL.scala 102:19]
  wire  m_604_io_x1; // @[MUL.scala 102:19]
  wire  m_604_io_x2; // @[MUL.scala 102:19]
  wire  m_604_io_x3; // @[MUL.scala 102:19]
  wire  m_604_io_s; // @[MUL.scala 102:19]
  wire  m_604_io_cout; // @[MUL.scala 102:19]
  wire  m_605_io_x1; // @[MUL.scala 102:19]
  wire  m_605_io_x2; // @[MUL.scala 102:19]
  wire  m_605_io_x3; // @[MUL.scala 102:19]
  wire  m_605_io_s; // @[MUL.scala 102:19]
  wire  m_605_io_cout; // @[MUL.scala 102:19]
  wire  m_606_io_x1; // @[MUL.scala 102:19]
  wire  m_606_io_x2; // @[MUL.scala 102:19]
  wire  m_606_io_x3; // @[MUL.scala 102:19]
  wire  m_606_io_s; // @[MUL.scala 102:19]
  wire  m_606_io_cout; // @[MUL.scala 102:19]
  wire  m_607_io_x1; // @[MUL.scala 102:19]
  wire  m_607_io_x2; // @[MUL.scala 102:19]
  wire  m_607_io_x3; // @[MUL.scala 102:19]
  wire  m_607_io_s; // @[MUL.scala 102:19]
  wire  m_607_io_cout; // @[MUL.scala 102:19]
  wire  m_608_io_x1; // @[MUL.scala 102:19]
  wire  m_608_io_x2; // @[MUL.scala 102:19]
  wire  m_608_io_x3; // @[MUL.scala 102:19]
  wire  m_608_io_s; // @[MUL.scala 102:19]
  wire  m_608_io_cout; // @[MUL.scala 102:19]
  wire  m_609_io_x1; // @[MUL.scala 102:19]
  wire  m_609_io_x2; // @[MUL.scala 102:19]
  wire  m_609_io_x3; // @[MUL.scala 102:19]
  wire  m_609_io_s; // @[MUL.scala 102:19]
  wire  m_609_io_cout; // @[MUL.scala 102:19]
  wire  m_610_io_x1; // @[MUL.scala 102:19]
  wire  m_610_io_x2; // @[MUL.scala 102:19]
  wire  m_610_io_x3; // @[MUL.scala 102:19]
  wire  m_610_io_s; // @[MUL.scala 102:19]
  wire  m_610_io_cout; // @[MUL.scala 102:19]
  wire  m_611_io_x1; // @[MUL.scala 102:19]
  wire  m_611_io_x2; // @[MUL.scala 102:19]
  wire  m_611_io_x3; // @[MUL.scala 102:19]
  wire  m_611_io_s; // @[MUL.scala 102:19]
  wire  m_611_io_cout; // @[MUL.scala 102:19]
  wire  m_612_io_x1; // @[MUL.scala 102:19]
  wire  m_612_io_x2; // @[MUL.scala 102:19]
  wire  m_612_io_x3; // @[MUL.scala 102:19]
  wire  m_612_io_s; // @[MUL.scala 102:19]
  wire  m_612_io_cout; // @[MUL.scala 102:19]
  wire  m_613_io_x1; // @[MUL.scala 102:19]
  wire  m_613_io_x2; // @[MUL.scala 102:19]
  wire  m_613_io_x3; // @[MUL.scala 102:19]
  wire  m_613_io_s; // @[MUL.scala 102:19]
  wire  m_613_io_cout; // @[MUL.scala 102:19]
  wire  m_614_io_x1; // @[MUL.scala 102:19]
  wire  m_614_io_x2; // @[MUL.scala 102:19]
  wire  m_614_io_x3; // @[MUL.scala 102:19]
  wire  m_614_io_s; // @[MUL.scala 102:19]
  wire  m_614_io_cout; // @[MUL.scala 102:19]
  wire  m_615_io_x1; // @[MUL.scala 102:19]
  wire  m_615_io_x2; // @[MUL.scala 102:19]
  wire  m_615_io_x3; // @[MUL.scala 102:19]
  wire  m_615_io_s; // @[MUL.scala 102:19]
  wire  m_615_io_cout; // @[MUL.scala 102:19]
  wire  m_616_io_x1; // @[MUL.scala 102:19]
  wire  m_616_io_x2; // @[MUL.scala 102:19]
  wire  m_616_io_x3; // @[MUL.scala 102:19]
  wire  m_616_io_s; // @[MUL.scala 102:19]
  wire  m_616_io_cout; // @[MUL.scala 102:19]
  wire  m_617_io_x1; // @[MUL.scala 102:19]
  wire  m_617_io_x2; // @[MUL.scala 102:19]
  wire  m_617_io_x3; // @[MUL.scala 102:19]
  wire  m_617_io_s; // @[MUL.scala 102:19]
  wire  m_617_io_cout; // @[MUL.scala 102:19]
  wire  m_618_io_x1; // @[MUL.scala 102:19]
  wire  m_618_io_x2; // @[MUL.scala 102:19]
  wire  m_618_io_x3; // @[MUL.scala 102:19]
  wire  m_618_io_s; // @[MUL.scala 102:19]
  wire  m_618_io_cout; // @[MUL.scala 102:19]
  wire  m_619_io_x1; // @[MUL.scala 102:19]
  wire  m_619_io_x2; // @[MUL.scala 102:19]
  wire  m_619_io_x3; // @[MUL.scala 102:19]
  wire  m_619_io_s; // @[MUL.scala 102:19]
  wire  m_619_io_cout; // @[MUL.scala 102:19]
  wire  m_620_io_x1; // @[MUL.scala 102:19]
  wire  m_620_io_x2; // @[MUL.scala 102:19]
  wire  m_620_io_x3; // @[MUL.scala 102:19]
  wire  m_620_io_s; // @[MUL.scala 102:19]
  wire  m_620_io_cout; // @[MUL.scala 102:19]
  wire  m_621_io_x1; // @[MUL.scala 102:19]
  wire  m_621_io_x2; // @[MUL.scala 102:19]
  wire  m_621_io_x3; // @[MUL.scala 102:19]
  wire  m_621_io_s; // @[MUL.scala 102:19]
  wire  m_621_io_cout; // @[MUL.scala 102:19]
  wire  m_622_io_x1; // @[MUL.scala 102:19]
  wire  m_622_io_x2; // @[MUL.scala 102:19]
  wire  m_622_io_x3; // @[MUL.scala 102:19]
  wire  m_622_io_s; // @[MUL.scala 102:19]
  wire  m_622_io_cout; // @[MUL.scala 102:19]
  wire  m_623_io_x1; // @[MUL.scala 102:19]
  wire  m_623_io_x2; // @[MUL.scala 102:19]
  wire  m_623_io_x3; // @[MUL.scala 102:19]
  wire  m_623_io_s; // @[MUL.scala 102:19]
  wire  m_623_io_cout; // @[MUL.scala 102:19]
  wire  m_624_io_x1; // @[MUL.scala 102:19]
  wire  m_624_io_x2; // @[MUL.scala 102:19]
  wire  m_624_io_x3; // @[MUL.scala 102:19]
  wire  m_624_io_s; // @[MUL.scala 102:19]
  wire  m_624_io_cout; // @[MUL.scala 102:19]
  wire  m_625_io_x1; // @[MUL.scala 102:19]
  wire  m_625_io_x2; // @[MUL.scala 102:19]
  wire  m_625_io_x3; // @[MUL.scala 102:19]
  wire  m_625_io_s; // @[MUL.scala 102:19]
  wire  m_625_io_cout; // @[MUL.scala 102:19]
  wire  m_626_io_in_0; // @[MUL.scala 124:19]
  wire  m_626_io_in_1; // @[MUL.scala 124:19]
  wire  m_626_io_out_0; // @[MUL.scala 124:19]
  wire  m_626_io_out_1; // @[MUL.scala 124:19]
  wire  m_627_io_x1; // @[MUL.scala 102:19]
  wire  m_627_io_x2; // @[MUL.scala 102:19]
  wire  m_627_io_x3; // @[MUL.scala 102:19]
  wire  m_627_io_s; // @[MUL.scala 102:19]
  wire  m_627_io_cout; // @[MUL.scala 102:19]
  wire  m_628_io_x1; // @[MUL.scala 102:19]
  wire  m_628_io_x2; // @[MUL.scala 102:19]
  wire  m_628_io_x3; // @[MUL.scala 102:19]
  wire  m_628_io_s; // @[MUL.scala 102:19]
  wire  m_628_io_cout; // @[MUL.scala 102:19]
  wire  m_629_io_x1; // @[MUL.scala 102:19]
  wire  m_629_io_x2; // @[MUL.scala 102:19]
  wire  m_629_io_x3; // @[MUL.scala 102:19]
  wire  m_629_io_s; // @[MUL.scala 102:19]
  wire  m_629_io_cout; // @[MUL.scala 102:19]
  wire  m_630_io_x1; // @[MUL.scala 102:19]
  wire  m_630_io_x2; // @[MUL.scala 102:19]
  wire  m_630_io_x3; // @[MUL.scala 102:19]
  wire  m_630_io_s; // @[MUL.scala 102:19]
  wire  m_630_io_cout; // @[MUL.scala 102:19]
  wire  m_631_io_x1; // @[MUL.scala 102:19]
  wire  m_631_io_x2; // @[MUL.scala 102:19]
  wire  m_631_io_x3; // @[MUL.scala 102:19]
  wire  m_631_io_s; // @[MUL.scala 102:19]
  wire  m_631_io_cout; // @[MUL.scala 102:19]
  wire  m_632_io_x1; // @[MUL.scala 102:19]
  wire  m_632_io_x2; // @[MUL.scala 102:19]
  wire  m_632_io_x3; // @[MUL.scala 102:19]
  wire  m_632_io_s; // @[MUL.scala 102:19]
  wire  m_632_io_cout; // @[MUL.scala 102:19]
  wire  m_633_io_x1; // @[MUL.scala 102:19]
  wire  m_633_io_x2; // @[MUL.scala 102:19]
  wire  m_633_io_x3; // @[MUL.scala 102:19]
  wire  m_633_io_s; // @[MUL.scala 102:19]
  wire  m_633_io_cout; // @[MUL.scala 102:19]
  wire  m_634_io_in_0; // @[MUL.scala 124:19]
  wire  m_634_io_in_1; // @[MUL.scala 124:19]
  wire  m_634_io_out_0; // @[MUL.scala 124:19]
  wire  m_634_io_out_1; // @[MUL.scala 124:19]
  wire  m_635_io_x1; // @[MUL.scala 102:19]
  wire  m_635_io_x2; // @[MUL.scala 102:19]
  wire  m_635_io_x3; // @[MUL.scala 102:19]
  wire  m_635_io_s; // @[MUL.scala 102:19]
  wire  m_635_io_cout; // @[MUL.scala 102:19]
  wire  m_636_io_x1; // @[MUL.scala 102:19]
  wire  m_636_io_x2; // @[MUL.scala 102:19]
  wire  m_636_io_x3; // @[MUL.scala 102:19]
  wire  m_636_io_s; // @[MUL.scala 102:19]
  wire  m_636_io_cout; // @[MUL.scala 102:19]
  wire  m_637_io_x1; // @[MUL.scala 102:19]
  wire  m_637_io_x2; // @[MUL.scala 102:19]
  wire  m_637_io_x3; // @[MUL.scala 102:19]
  wire  m_637_io_s; // @[MUL.scala 102:19]
  wire  m_637_io_cout; // @[MUL.scala 102:19]
  wire  m_638_io_x1; // @[MUL.scala 102:19]
  wire  m_638_io_x2; // @[MUL.scala 102:19]
  wire  m_638_io_x3; // @[MUL.scala 102:19]
  wire  m_638_io_s; // @[MUL.scala 102:19]
  wire  m_638_io_cout; // @[MUL.scala 102:19]
  wire  m_639_io_x1; // @[MUL.scala 102:19]
  wire  m_639_io_x2; // @[MUL.scala 102:19]
  wire  m_639_io_x3; // @[MUL.scala 102:19]
  wire  m_639_io_s; // @[MUL.scala 102:19]
  wire  m_639_io_cout; // @[MUL.scala 102:19]
  wire  m_640_io_x1; // @[MUL.scala 102:19]
  wire  m_640_io_x2; // @[MUL.scala 102:19]
  wire  m_640_io_x3; // @[MUL.scala 102:19]
  wire  m_640_io_s; // @[MUL.scala 102:19]
  wire  m_640_io_cout; // @[MUL.scala 102:19]
  wire  m_641_io_x1; // @[MUL.scala 102:19]
  wire  m_641_io_x2; // @[MUL.scala 102:19]
  wire  m_641_io_x3; // @[MUL.scala 102:19]
  wire  m_641_io_s; // @[MUL.scala 102:19]
  wire  m_641_io_cout; // @[MUL.scala 102:19]
  wire  m_642_io_x1; // @[MUL.scala 102:19]
  wire  m_642_io_x2; // @[MUL.scala 102:19]
  wire  m_642_io_x3; // @[MUL.scala 102:19]
  wire  m_642_io_s; // @[MUL.scala 102:19]
  wire  m_642_io_cout; // @[MUL.scala 102:19]
  wire  m_643_io_x1; // @[MUL.scala 102:19]
  wire  m_643_io_x2; // @[MUL.scala 102:19]
  wire  m_643_io_x3; // @[MUL.scala 102:19]
  wire  m_643_io_s; // @[MUL.scala 102:19]
  wire  m_643_io_cout; // @[MUL.scala 102:19]
  wire  m_644_io_x1; // @[MUL.scala 102:19]
  wire  m_644_io_x2; // @[MUL.scala 102:19]
  wire  m_644_io_x3; // @[MUL.scala 102:19]
  wire  m_644_io_s; // @[MUL.scala 102:19]
  wire  m_644_io_cout; // @[MUL.scala 102:19]
  wire  m_645_io_x1; // @[MUL.scala 102:19]
  wire  m_645_io_x2; // @[MUL.scala 102:19]
  wire  m_645_io_x3; // @[MUL.scala 102:19]
  wire  m_645_io_s; // @[MUL.scala 102:19]
  wire  m_645_io_cout; // @[MUL.scala 102:19]
  wire  m_646_io_x1; // @[MUL.scala 102:19]
  wire  m_646_io_x2; // @[MUL.scala 102:19]
  wire  m_646_io_x3; // @[MUL.scala 102:19]
  wire  m_646_io_s; // @[MUL.scala 102:19]
  wire  m_646_io_cout; // @[MUL.scala 102:19]
  wire  m_647_io_x1; // @[MUL.scala 102:19]
  wire  m_647_io_x2; // @[MUL.scala 102:19]
  wire  m_647_io_x3; // @[MUL.scala 102:19]
  wire  m_647_io_s; // @[MUL.scala 102:19]
  wire  m_647_io_cout; // @[MUL.scala 102:19]
  wire  m_648_io_x1; // @[MUL.scala 102:19]
  wire  m_648_io_x2; // @[MUL.scala 102:19]
  wire  m_648_io_x3; // @[MUL.scala 102:19]
  wire  m_648_io_s; // @[MUL.scala 102:19]
  wire  m_648_io_cout; // @[MUL.scala 102:19]
  wire  m_649_io_x1; // @[MUL.scala 102:19]
  wire  m_649_io_x2; // @[MUL.scala 102:19]
  wire  m_649_io_x3; // @[MUL.scala 102:19]
  wire  m_649_io_s; // @[MUL.scala 102:19]
  wire  m_649_io_cout; // @[MUL.scala 102:19]
  wire  m_650_io_x1; // @[MUL.scala 102:19]
  wire  m_650_io_x2; // @[MUL.scala 102:19]
  wire  m_650_io_x3; // @[MUL.scala 102:19]
  wire  m_650_io_s; // @[MUL.scala 102:19]
  wire  m_650_io_cout; // @[MUL.scala 102:19]
  wire  m_651_io_x1; // @[MUL.scala 102:19]
  wire  m_651_io_x2; // @[MUL.scala 102:19]
  wire  m_651_io_x3; // @[MUL.scala 102:19]
  wire  m_651_io_s; // @[MUL.scala 102:19]
  wire  m_651_io_cout; // @[MUL.scala 102:19]
  wire  m_652_io_x1; // @[MUL.scala 102:19]
  wire  m_652_io_x2; // @[MUL.scala 102:19]
  wire  m_652_io_x3; // @[MUL.scala 102:19]
  wire  m_652_io_s; // @[MUL.scala 102:19]
  wire  m_652_io_cout; // @[MUL.scala 102:19]
  wire  m_653_io_x1; // @[MUL.scala 102:19]
  wire  m_653_io_x2; // @[MUL.scala 102:19]
  wire  m_653_io_x3; // @[MUL.scala 102:19]
  wire  m_653_io_s; // @[MUL.scala 102:19]
  wire  m_653_io_cout; // @[MUL.scala 102:19]
  wire  m_654_io_x1; // @[MUL.scala 102:19]
  wire  m_654_io_x2; // @[MUL.scala 102:19]
  wire  m_654_io_x3; // @[MUL.scala 102:19]
  wire  m_654_io_s; // @[MUL.scala 102:19]
  wire  m_654_io_cout; // @[MUL.scala 102:19]
  wire  m_655_io_x1; // @[MUL.scala 102:19]
  wire  m_655_io_x2; // @[MUL.scala 102:19]
  wire  m_655_io_x3; // @[MUL.scala 102:19]
  wire  m_655_io_s; // @[MUL.scala 102:19]
  wire  m_655_io_cout; // @[MUL.scala 102:19]
  wire  m_656_io_x1; // @[MUL.scala 102:19]
  wire  m_656_io_x2; // @[MUL.scala 102:19]
  wire  m_656_io_x3; // @[MUL.scala 102:19]
  wire  m_656_io_s; // @[MUL.scala 102:19]
  wire  m_656_io_cout; // @[MUL.scala 102:19]
  wire  m_657_io_x1; // @[MUL.scala 102:19]
  wire  m_657_io_x2; // @[MUL.scala 102:19]
  wire  m_657_io_x3; // @[MUL.scala 102:19]
  wire  m_657_io_s; // @[MUL.scala 102:19]
  wire  m_657_io_cout; // @[MUL.scala 102:19]
  wire  m_658_io_x1; // @[MUL.scala 102:19]
  wire  m_658_io_x2; // @[MUL.scala 102:19]
  wire  m_658_io_x3; // @[MUL.scala 102:19]
  wire  m_658_io_s; // @[MUL.scala 102:19]
  wire  m_658_io_cout; // @[MUL.scala 102:19]
  wire  m_659_io_x1; // @[MUL.scala 102:19]
  wire  m_659_io_x2; // @[MUL.scala 102:19]
  wire  m_659_io_x3; // @[MUL.scala 102:19]
  wire  m_659_io_s; // @[MUL.scala 102:19]
  wire  m_659_io_cout; // @[MUL.scala 102:19]
  wire  m_660_io_x1; // @[MUL.scala 102:19]
  wire  m_660_io_x2; // @[MUL.scala 102:19]
  wire  m_660_io_x3; // @[MUL.scala 102:19]
  wire  m_660_io_s; // @[MUL.scala 102:19]
  wire  m_660_io_cout; // @[MUL.scala 102:19]
  wire  m_661_io_x1; // @[MUL.scala 102:19]
  wire  m_661_io_x2; // @[MUL.scala 102:19]
  wire  m_661_io_x3; // @[MUL.scala 102:19]
  wire  m_661_io_s; // @[MUL.scala 102:19]
  wire  m_661_io_cout; // @[MUL.scala 102:19]
  wire  m_662_io_x1; // @[MUL.scala 102:19]
  wire  m_662_io_x2; // @[MUL.scala 102:19]
  wire  m_662_io_x3; // @[MUL.scala 102:19]
  wire  m_662_io_s; // @[MUL.scala 102:19]
  wire  m_662_io_cout; // @[MUL.scala 102:19]
  wire  m_663_io_x1; // @[MUL.scala 102:19]
  wire  m_663_io_x2; // @[MUL.scala 102:19]
  wire  m_663_io_x3; // @[MUL.scala 102:19]
  wire  m_663_io_s; // @[MUL.scala 102:19]
  wire  m_663_io_cout; // @[MUL.scala 102:19]
  wire  m_664_io_x1; // @[MUL.scala 102:19]
  wire  m_664_io_x2; // @[MUL.scala 102:19]
  wire  m_664_io_x3; // @[MUL.scala 102:19]
  wire  m_664_io_s; // @[MUL.scala 102:19]
  wire  m_664_io_cout; // @[MUL.scala 102:19]
  wire  m_665_io_x1; // @[MUL.scala 102:19]
  wire  m_665_io_x2; // @[MUL.scala 102:19]
  wire  m_665_io_x3; // @[MUL.scala 102:19]
  wire  m_665_io_s; // @[MUL.scala 102:19]
  wire  m_665_io_cout; // @[MUL.scala 102:19]
  wire  m_666_io_x1; // @[MUL.scala 102:19]
  wire  m_666_io_x2; // @[MUL.scala 102:19]
  wire  m_666_io_x3; // @[MUL.scala 102:19]
  wire  m_666_io_s; // @[MUL.scala 102:19]
  wire  m_666_io_cout; // @[MUL.scala 102:19]
  wire  m_667_io_x1; // @[MUL.scala 102:19]
  wire  m_667_io_x2; // @[MUL.scala 102:19]
  wire  m_667_io_x3; // @[MUL.scala 102:19]
  wire  m_667_io_s; // @[MUL.scala 102:19]
  wire  m_667_io_cout; // @[MUL.scala 102:19]
  wire  m_668_io_x1; // @[MUL.scala 102:19]
  wire  m_668_io_x2; // @[MUL.scala 102:19]
  wire  m_668_io_x3; // @[MUL.scala 102:19]
  wire  m_668_io_s; // @[MUL.scala 102:19]
  wire  m_668_io_cout; // @[MUL.scala 102:19]
  wire  m_669_io_in_0; // @[MUL.scala 124:19]
  wire  m_669_io_in_1; // @[MUL.scala 124:19]
  wire  m_669_io_out_0; // @[MUL.scala 124:19]
  wire  m_669_io_out_1; // @[MUL.scala 124:19]
  wire  m_670_io_x1; // @[MUL.scala 102:19]
  wire  m_670_io_x2; // @[MUL.scala 102:19]
  wire  m_670_io_x3; // @[MUL.scala 102:19]
  wire  m_670_io_s; // @[MUL.scala 102:19]
  wire  m_670_io_cout; // @[MUL.scala 102:19]
  wire  m_671_io_x1; // @[MUL.scala 102:19]
  wire  m_671_io_x2; // @[MUL.scala 102:19]
  wire  m_671_io_x3; // @[MUL.scala 102:19]
  wire  m_671_io_s; // @[MUL.scala 102:19]
  wire  m_671_io_cout; // @[MUL.scala 102:19]
  wire  m_672_io_x1; // @[MUL.scala 102:19]
  wire  m_672_io_x2; // @[MUL.scala 102:19]
  wire  m_672_io_x3; // @[MUL.scala 102:19]
  wire  m_672_io_s; // @[MUL.scala 102:19]
  wire  m_672_io_cout; // @[MUL.scala 102:19]
  wire  m_673_io_x1; // @[MUL.scala 102:19]
  wire  m_673_io_x2; // @[MUL.scala 102:19]
  wire  m_673_io_x3; // @[MUL.scala 102:19]
  wire  m_673_io_s; // @[MUL.scala 102:19]
  wire  m_673_io_cout; // @[MUL.scala 102:19]
  wire  m_674_io_x1; // @[MUL.scala 102:19]
  wire  m_674_io_x2; // @[MUL.scala 102:19]
  wire  m_674_io_x3; // @[MUL.scala 102:19]
  wire  m_674_io_s; // @[MUL.scala 102:19]
  wire  m_674_io_cout; // @[MUL.scala 102:19]
  wire  m_675_io_x1; // @[MUL.scala 102:19]
  wire  m_675_io_x2; // @[MUL.scala 102:19]
  wire  m_675_io_x3; // @[MUL.scala 102:19]
  wire  m_675_io_s; // @[MUL.scala 102:19]
  wire  m_675_io_cout; // @[MUL.scala 102:19]
  wire  m_676_io_in_0; // @[MUL.scala 124:19]
  wire  m_676_io_in_1; // @[MUL.scala 124:19]
  wire  m_676_io_out_0; // @[MUL.scala 124:19]
  wire  m_676_io_out_1; // @[MUL.scala 124:19]
  wire  m_677_io_x1; // @[MUL.scala 102:19]
  wire  m_677_io_x2; // @[MUL.scala 102:19]
  wire  m_677_io_x3; // @[MUL.scala 102:19]
  wire  m_677_io_s; // @[MUL.scala 102:19]
  wire  m_677_io_cout; // @[MUL.scala 102:19]
  wire  m_678_io_x1; // @[MUL.scala 102:19]
  wire  m_678_io_x2; // @[MUL.scala 102:19]
  wire  m_678_io_x3; // @[MUL.scala 102:19]
  wire  m_678_io_s; // @[MUL.scala 102:19]
  wire  m_678_io_cout; // @[MUL.scala 102:19]
  wire  m_679_io_x1; // @[MUL.scala 102:19]
  wire  m_679_io_x2; // @[MUL.scala 102:19]
  wire  m_679_io_x3; // @[MUL.scala 102:19]
  wire  m_679_io_s; // @[MUL.scala 102:19]
  wire  m_679_io_cout; // @[MUL.scala 102:19]
  wire  m_680_io_x1; // @[MUL.scala 102:19]
  wire  m_680_io_x2; // @[MUL.scala 102:19]
  wire  m_680_io_x3; // @[MUL.scala 102:19]
  wire  m_680_io_s; // @[MUL.scala 102:19]
  wire  m_680_io_cout; // @[MUL.scala 102:19]
  wire  m_681_io_x1; // @[MUL.scala 102:19]
  wire  m_681_io_x2; // @[MUL.scala 102:19]
  wire  m_681_io_x3; // @[MUL.scala 102:19]
  wire  m_681_io_s; // @[MUL.scala 102:19]
  wire  m_681_io_cout; // @[MUL.scala 102:19]
  wire  m_682_io_x1; // @[MUL.scala 102:19]
  wire  m_682_io_x2; // @[MUL.scala 102:19]
  wire  m_682_io_x3; // @[MUL.scala 102:19]
  wire  m_682_io_s; // @[MUL.scala 102:19]
  wire  m_682_io_cout; // @[MUL.scala 102:19]
  wire  m_683_io_x1; // @[MUL.scala 102:19]
  wire  m_683_io_x2; // @[MUL.scala 102:19]
  wire  m_683_io_x3; // @[MUL.scala 102:19]
  wire  m_683_io_s; // @[MUL.scala 102:19]
  wire  m_683_io_cout; // @[MUL.scala 102:19]
  wire  m_684_io_x1; // @[MUL.scala 102:19]
  wire  m_684_io_x2; // @[MUL.scala 102:19]
  wire  m_684_io_x3; // @[MUL.scala 102:19]
  wire  m_684_io_s; // @[MUL.scala 102:19]
  wire  m_684_io_cout; // @[MUL.scala 102:19]
  wire  m_685_io_x1; // @[MUL.scala 102:19]
  wire  m_685_io_x2; // @[MUL.scala 102:19]
  wire  m_685_io_x3; // @[MUL.scala 102:19]
  wire  m_685_io_s; // @[MUL.scala 102:19]
  wire  m_685_io_cout; // @[MUL.scala 102:19]
  wire  m_686_io_x1; // @[MUL.scala 102:19]
  wire  m_686_io_x2; // @[MUL.scala 102:19]
  wire  m_686_io_x3; // @[MUL.scala 102:19]
  wire  m_686_io_s; // @[MUL.scala 102:19]
  wire  m_686_io_cout; // @[MUL.scala 102:19]
  wire  m_687_io_x1; // @[MUL.scala 102:19]
  wire  m_687_io_x2; // @[MUL.scala 102:19]
  wire  m_687_io_x3; // @[MUL.scala 102:19]
  wire  m_687_io_s; // @[MUL.scala 102:19]
  wire  m_687_io_cout; // @[MUL.scala 102:19]
  wire  m_688_io_x1; // @[MUL.scala 102:19]
  wire  m_688_io_x2; // @[MUL.scala 102:19]
  wire  m_688_io_x3; // @[MUL.scala 102:19]
  wire  m_688_io_s; // @[MUL.scala 102:19]
  wire  m_688_io_cout; // @[MUL.scala 102:19]
  wire  m_689_io_x1; // @[MUL.scala 102:19]
  wire  m_689_io_x2; // @[MUL.scala 102:19]
  wire  m_689_io_x3; // @[MUL.scala 102:19]
  wire  m_689_io_s; // @[MUL.scala 102:19]
  wire  m_689_io_cout; // @[MUL.scala 102:19]
  wire  m_690_io_x1; // @[MUL.scala 102:19]
  wire  m_690_io_x2; // @[MUL.scala 102:19]
  wire  m_690_io_x3; // @[MUL.scala 102:19]
  wire  m_690_io_s; // @[MUL.scala 102:19]
  wire  m_690_io_cout; // @[MUL.scala 102:19]
  wire  m_691_io_x1; // @[MUL.scala 102:19]
  wire  m_691_io_x2; // @[MUL.scala 102:19]
  wire  m_691_io_x3; // @[MUL.scala 102:19]
  wire  m_691_io_s; // @[MUL.scala 102:19]
  wire  m_691_io_cout; // @[MUL.scala 102:19]
  wire  m_692_io_x1; // @[MUL.scala 102:19]
  wire  m_692_io_x2; // @[MUL.scala 102:19]
  wire  m_692_io_x3; // @[MUL.scala 102:19]
  wire  m_692_io_s; // @[MUL.scala 102:19]
  wire  m_692_io_cout; // @[MUL.scala 102:19]
  wire  m_693_io_x1; // @[MUL.scala 102:19]
  wire  m_693_io_x2; // @[MUL.scala 102:19]
  wire  m_693_io_x3; // @[MUL.scala 102:19]
  wire  m_693_io_s; // @[MUL.scala 102:19]
  wire  m_693_io_cout; // @[MUL.scala 102:19]
  wire  m_694_io_x1; // @[MUL.scala 102:19]
  wire  m_694_io_x2; // @[MUL.scala 102:19]
  wire  m_694_io_x3; // @[MUL.scala 102:19]
  wire  m_694_io_s; // @[MUL.scala 102:19]
  wire  m_694_io_cout; // @[MUL.scala 102:19]
  wire  m_695_io_x1; // @[MUL.scala 102:19]
  wire  m_695_io_x2; // @[MUL.scala 102:19]
  wire  m_695_io_x3; // @[MUL.scala 102:19]
  wire  m_695_io_s; // @[MUL.scala 102:19]
  wire  m_695_io_cout; // @[MUL.scala 102:19]
  wire  m_696_io_x1; // @[MUL.scala 102:19]
  wire  m_696_io_x2; // @[MUL.scala 102:19]
  wire  m_696_io_x3; // @[MUL.scala 102:19]
  wire  m_696_io_s; // @[MUL.scala 102:19]
  wire  m_696_io_cout; // @[MUL.scala 102:19]
  wire  m_697_io_x1; // @[MUL.scala 102:19]
  wire  m_697_io_x2; // @[MUL.scala 102:19]
  wire  m_697_io_x3; // @[MUL.scala 102:19]
  wire  m_697_io_s; // @[MUL.scala 102:19]
  wire  m_697_io_cout; // @[MUL.scala 102:19]
  wire  m_698_io_x1; // @[MUL.scala 102:19]
  wire  m_698_io_x2; // @[MUL.scala 102:19]
  wire  m_698_io_x3; // @[MUL.scala 102:19]
  wire  m_698_io_s; // @[MUL.scala 102:19]
  wire  m_698_io_cout; // @[MUL.scala 102:19]
  wire  m_699_io_x1; // @[MUL.scala 102:19]
  wire  m_699_io_x2; // @[MUL.scala 102:19]
  wire  m_699_io_x3; // @[MUL.scala 102:19]
  wire  m_699_io_s; // @[MUL.scala 102:19]
  wire  m_699_io_cout; // @[MUL.scala 102:19]
  wire  m_700_io_x1; // @[MUL.scala 102:19]
  wire  m_700_io_x2; // @[MUL.scala 102:19]
  wire  m_700_io_x3; // @[MUL.scala 102:19]
  wire  m_700_io_s; // @[MUL.scala 102:19]
  wire  m_700_io_cout; // @[MUL.scala 102:19]
  wire  m_701_io_x1; // @[MUL.scala 102:19]
  wire  m_701_io_x2; // @[MUL.scala 102:19]
  wire  m_701_io_x3; // @[MUL.scala 102:19]
  wire  m_701_io_s; // @[MUL.scala 102:19]
  wire  m_701_io_cout; // @[MUL.scala 102:19]
  wire  m_702_io_x1; // @[MUL.scala 102:19]
  wire  m_702_io_x2; // @[MUL.scala 102:19]
  wire  m_702_io_x3; // @[MUL.scala 102:19]
  wire  m_702_io_s; // @[MUL.scala 102:19]
  wire  m_702_io_cout; // @[MUL.scala 102:19]
  wire  m_703_io_x1; // @[MUL.scala 102:19]
  wire  m_703_io_x2; // @[MUL.scala 102:19]
  wire  m_703_io_x3; // @[MUL.scala 102:19]
  wire  m_703_io_s; // @[MUL.scala 102:19]
  wire  m_703_io_cout; // @[MUL.scala 102:19]
  wire  m_704_io_x1; // @[MUL.scala 102:19]
  wire  m_704_io_x2; // @[MUL.scala 102:19]
  wire  m_704_io_x3; // @[MUL.scala 102:19]
  wire  m_704_io_s; // @[MUL.scala 102:19]
  wire  m_704_io_cout; // @[MUL.scala 102:19]
  wire  m_705_io_x1; // @[MUL.scala 102:19]
  wire  m_705_io_x2; // @[MUL.scala 102:19]
  wire  m_705_io_x3; // @[MUL.scala 102:19]
  wire  m_705_io_s; // @[MUL.scala 102:19]
  wire  m_705_io_cout; // @[MUL.scala 102:19]
  wire  m_706_io_in_0; // @[MUL.scala 124:19]
  wire  m_706_io_in_1; // @[MUL.scala 124:19]
  wire  m_706_io_out_0; // @[MUL.scala 124:19]
  wire  m_706_io_out_1; // @[MUL.scala 124:19]
  wire  m_707_io_x1; // @[MUL.scala 102:19]
  wire  m_707_io_x2; // @[MUL.scala 102:19]
  wire  m_707_io_x3; // @[MUL.scala 102:19]
  wire  m_707_io_s; // @[MUL.scala 102:19]
  wire  m_707_io_cout; // @[MUL.scala 102:19]
  wire  m_708_io_x1; // @[MUL.scala 102:19]
  wire  m_708_io_x2; // @[MUL.scala 102:19]
  wire  m_708_io_x3; // @[MUL.scala 102:19]
  wire  m_708_io_s; // @[MUL.scala 102:19]
  wire  m_708_io_cout; // @[MUL.scala 102:19]
  wire  m_709_io_x1; // @[MUL.scala 102:19]
  wire  m_709_io_x2; // @[MUL.scala 102:19]
  wire  m_709_io_x3; // @[MUL.scala 102:19]
  wire  m_709_io_s; // @[MUL.scala 102:19]
  wire  m_709_io_cout; // @[MUL.scala 102:19]
  wire  m_710_io_x1; // @[MUL.scala 102:19]
  wire  m_710_io_x2; // @[MUL.scala 102:19]
  wire  m_710_io_x3; // @[MUL.scala 102:19]
  wire  m_710_io_s; // @[MUL.scala 102:19]
  wire  m_710_io_cout; // @[MUL.scala 102:19]
  wire  m_711_io_x1; // @[MUL.scala 102:19]
  wire  m_711_io_x2; // @[MUL.scala 102:19]
  wire  m_711_io_x3; // @[MUL.scala 102:19]
  wire  m_711_io_s; // @[MUL.scala 102:19]
  wire  m_711_io_cout; // @[MUL.scala 102:19]
  wire  m_712_io_in_0; // @[MUL.scala 124:19]
  wire  m_712_io_in_1; // @[MUL.scala 124:19]
  wire  m_712_io_out_0; // @[MUL.scala 124:19]
  wire  m_712_io_out_1; // @[MUL.scala 124:19]
  wire  m_713_io_x1; // @[MUL.scala 102:19]
  wire  m_713_io_x2; // @[MUL.scala 102:19]
  wire  m_713_io_x3; // @[MUL.scala 102:19]
  wire  m_713_io_s; // @[MUL.scala 102:19]
  wire  m_713_io_cout; // @[MUL.scala 102:19]
  wire  m_714_io_x1; // @[MUL.scala 102:19]
  wire  m_714_io_x2; // @[MUL.scala 102:19]
  wire  m_714_io_x3; // @[MUL.scala 102:19]
  wire  m_714_io_s; // @[MUL.scala 102:19]
  wire  m_714_io_cout; // @[MUL.scala 102:19]
  wire  m_715_io_x1; // @[MUL.scala 102:19]
  wire  m_715_io_x2; // @[MUL.scala 102:19]
  wire  m_715_io_x3; // @[MUL.scala 102:19]
  wire  m_715_io_s; // @[MUL.scala 102:19]
  wire  m_715_io_cout; // @[MUL.scala 102:19]
  wire  m_716_io_x1; // @[MUL.scala 102:19]
  wire  m_716_io_x2; // @[MUL.scala 102:19]
  wire  m_716_io_x3; // @[MUL.scala 102:19]
  wire  m_716_io_s; // @[MUL.scala 102:19]
  wire  m_716_io_cout; // @[MUL.scala 102:19]
  wire  m_717_io_x1; // @[MUL.scala 102:19]
  wire  m_717_io_x2; // @[MUL.scala 102:19]
  wire  m_717_io_x3; // @[MUL.scala 102:19]
  wire  m_717_io_s; // @[MUL.scala 102:19]
  wire  m_717_io_cout; // @[MUL.scala 102:19]
  wire  m_718_io_x1; // @[MUL.scala 102:19]
  wire  m_718_io_x2; // @[MUL.scala 102:19]
  wire  m_718_io_x3; // @[MUL.scala 102:19]
  wire  m_718_io_s; // @[MUL.scala 102:19]
  wire  m_718_io_cout; // @[MUL.scala 102:19]
  wire  m_719_io_x1; // @[MUL.scala 102:19]
  wire  m_719_io_x2; // @[MUL.scala 102:19]
  wire  m_719_io_x3; // @[MUL.scala 102:19]
  wire  m_719_io_s; // @[MUL.scala 102:19]
  wire  m_719_io_cout; // @[MUL.scala 102:19]
  wire  m_720_io_x1; // @[MUL.scala 102:19]
  wire  m_720_io_x2; // @[MUL.scala 102:19]
  wire  m_720_io_x3; // @[MUL.scala 102:19]
  wire  m_720_io_s; // @[MUL.scala 102:19]
  wire  m_720_io_cout; // @[MUL.scala 102:19]
  wire  m_721_io_x1; // @[MUL.scala 102:19]
  wire  m_721_io_x2; // @[MUL.scala 102:19]
  wire  m_721_io_x3; // @[MUL.scala 102:19]
  wire  m_721_io_s; // @[MUL.scala 102:19]
  wire  m_721_io_cout; // @[MUL.scala 102:19]
  wire  m_722_io_x1; // @[MUL.scala 102:19]
  wire  m_722_io_x2; // @[MUL.scala 102:19]
  wire  m_722_io_x3; // @[MUL.scala 102:19]
  wire  m_722_io_s; // @[MUL.scala 102:19]
  wire  m_722_io_cout; // @[MUL.scala 102:19]
  wire  m_723_io_x1; // @[MUL.scala 102:19]
  wire  m_723_io_x2; // @[MUL.scala 102:19]
  wire  m_723_io_x3; // @[MUL.scala 102:19]
  wire  m_723_io_s; // @[MUL.scala 102:19]
  wire  m_723_io_cout; // @[MUL.scala 102:19]
  wire  m_724_io_x1; // @[MUL.scala 102:19]
  wire  m_724_io_x2; // @[MUL.scala 102:19]
  wire  m_724_io_x3; // @[MUL.scala 102:19]
  wire  m_724_io_s; // @[MUL.scala 102:19]
  wire  m_724_io_cout; // @[MUL.scala 102:19]
  wire  m_725_io_x1; // @[MUL.scala 102:19]
  wire  m_725_io_x2; // @[MUL.scala 102:19]
  wire  m_725_io_x3; // @[MUL.scala 102:19]
  wire  m_725_io_s; // @[MUL.scala 102:19]
  wire  m_725_io_cout; // @[MUL.scala 102:19]
  wire  m_726_io_x1; // @[MUL.scala 102:19]
  wire  m_726_io_x2; // @[MUL.scala 102:19]
  wire  m_726_io_x3; // @[MUL.scala 102:19]
  wire  m_726_io_s; // @[MUL.scala 102:19]
  wire  m_726_io_cout; // @[MUL.scala 102:19]
  wire  m_727_io_x1; // @[MUL.scala 102:19]
  wire  m_727_io_x2; // @[MUL.scala 102:19]
  wire  m_727_io_x3; // @[MUL.scala 102:19]
  wire  m_727_io_s; // @[MUL.scala 102:19]
  wire  m_727_io_cout; // @[MUL.scala 102:19]
  wire  m_728_io_x1; // @[MUL.scala 102:19]
  wire  m_728_io_x2; // @[MUL.scala 102:19]
  wire  m_728_io_x3; // @[MUL.scala 102:19]
  wire  m_728_io_s; // @[MUL.scala 102:19]
  wire  m_728_io_cout; // @[MUL.scala 102:19]
  wire  m_729_io_x1; // @[MUL.scala 102:19]
  wire  m_729_io_x2; // @[MUL.scala 102:19]
  wire  m_729_io_x3; // @[MUL.scala 102:19]
  wire  m_729_io_s; // @[MUL.scala 102:19]
  wire  m_729_io_cout; // @[MUL.scala 102:19]
  wire  m_730_io_x1; // @[MUL.scala 102:19]
  wire  m_730_io_x2; // @[MUL.scala 102:19]
  wire  m_730_io_x3; // @[MUL.scala 102:19]
  wire  m_730_io_s; // @[MUL.scala 102:19]
  wire  m_730_io_cout; // @[MUL.scala 102:19]
  wire  m_731_io_x1; // @[MUL.scala 102:19]
  wire  m_731_io_x2; // @[MUL.scala 102:19]
  wire  m_731_io_x3; // @[MUL.scala 102:19]
  wire  m_731_io_s; // @[MUL.scala 102:19]
  wire  m_731_io_cout; // @[MUL.scala 102:19]
  wire  m_732_io_x1; // @[MUL.scala 102:19]
  wire  m_732_io_x2; // @[MUL.scala 102:19]
  wire  m_732_io_x3; // @[MUL.scala 102:19]
  wire  m_732_io_s; // @[MUL.scala 102:19]
  wire  m_732_io_cout; // @[MUL.scala 102:19]
  wire  m_733_io_x1; // @[MUL.scala 102:19]
  wire  m_733_io_x2; // @[MUL.scala 102:19]
  wire  m_733_io_x3; // @[MUL.scala 102:19]
  wire  m_733_io_s; // @[MUL.scala 102:19]
  wire  m_733_io_cout; // @[MUL.scala 102:19]
  wire  m_734_io_x1; // @[MUL.scala 102:19]
  wire  m_734_io_x2; // @[MUL.scala 102:19]
  wire  m_734_io_x3; // @[MUL.scala 102:19]
  wire  m_734_io_s; // @[MUL.scala 102:19]
  wire  m_734_io_cout; // @[MUL.scala 102:19]
  wire  m_735_io_x1; // @[MUL.scala 102:19]
  wire  m_735_io_x2; // @[MUL.scala 102:19]
  wire  m_735_io_x3; // @[MUL.scala 102:19]
  wire  m_735_io_s; // @[MUL.scala 102:19]
  wire  m_735_io_cout; // @[MUL.scala 102:19]
  wire  m_736_io_x1; // @[MUL.scala 102:19]
  wire  m_736_io_x2; // @[MUL.scala 102:19]
  wire  m_736_io_x3; // @[MUL.scala 102:19]
  wire  m_736_io_s; // @[MUL.scala 102:19]
  wire  m_736_io_cout; // @[MUL.scala 102:19]
  wire  m_737_io_in_0; // @[MUL.scala 124:19]
  wire  m_737_io_in_1; // @[MUL.scala 124:19]
  wire  m_737_io_out_0; // @[MUL.scala 124:19]
  wire  m_737_io_out_1; // @[MUL.scala 124:19]
  wire  m_738_io_x1; // @[MUL.scala 102:19]
  wire  m_738_io_x2; // @[MUL.scala 102:19]
  wire  m_738_io_x3; // @[MUL.scala 102:19]
  wire  m_738_io_s; // @[MUL.scala 102:19]
  wire  m_738_io_cout; // @[MUL.scala 102:19]
  wire  m_739_io_x1; // @[MUL.scala 102:19]
  wire  m_739_io_x2; // @[MUL.scala 102:19]
  wire  m_739_io_x3; // @[MUL.scala 102:19]
  wire  m_739_io_s; // @[MUL.scala 102:19]
  wire  m_739_io_cout; // @[MUL.scala 102:19]
  wire  m_740_io_x1; // @[MUL.scala 102:19]
  wire  m_740_io_x2; // @[MUL.scala 102:19]
  wire  m_740_io_x3; // @[MUL.scala 102:19]
  wire  m_740_io_s; // @[MUL.scala 102:19]
  wire  m_740_io_cout; // @[MUL.scala 102:19]
  wire  m_741_io_x1; // @[MUL.scala 102:19]
  wire  m_741_io_x2; // @[MUL.scala 102:19]
  wire  m_741_io_x3; // @[MUL.scala 102:19]
  wire  m_741_io_s; // @[MUL.scala 102:19]
  wire  m_741_io_cout; // @[MUL.scala 102:19]
  wire  m_742_io_in_0; // @[MUL.scala 124:19]
  wire  m_742_io_in_1; // @[MUL.scala 124:19]
  wire  m_742_io_out_0; // @[MUL.scala 124:19]
  wire  m_742_io_out_1; // @[MUL.scala 124:19]
  wire  m_743_io_x1; // @[MUL.scala 102:19]
  wire  m_743_io_x2; // @[MUL.scala 102:19]
  wire  m_743_io_x3; // @[MUL.scala 102:19]
  wire  m_743_io_s; // @[MUL.scala 102:19]
  wire  m_743_io_cout; // @[MUL.scala 102:19]
  wire  m_744_io_x1; // @[MUL.scala 102:19]
  wire  m_744_io_x2; // @[MUL.scala 102:19]
  wire  m_744_io_x3; // @[MUL.scala 102:19]
  wire  m_744_io_s; // @[MUL.scala 102:19]
  wire  m_744_io_cout; // @[MUL.scala 102:19]
  wire  m_745_io_x1; // @[MUL.scala 102:19]
  wire  m_745_io_x2; // @[MUL.scala 102:19]
  wire  m_745_io_x3; // @[MUL.scala 102:19]
  wire  m_745_io_s; // @[MUL.scala 102:19]
  wire  m_745_io_cout; // @[MUL.scala 102:19]
  wire  m_746_io_x1; // @[MUL.scala 102:19]
  wire  m_746_io_x2; // @[MUL.scala 102:19]
  wire  m_746_io_x3; // @[MUL.scala 102:19]
  wire  m_746_io_s; // @[MUL.scala 102:19]
  wire  m_746_io_cout; // @[MUL.scala 102:19]
  wire  m_747_io_x1; // @[MUL.scala 102:19]
  wire  m_747_io_x2; // @[MUL.scala 102:19]
  wire  m_747_io_x3; // @[MUL.scala 102:19]
  wire  m_747_io_s; // @[MUL.scala 102:19]
  wire  m_747_io_cout; // @[MUL.scala 102:19]
  wire  m_748_io_x1; // @[MUL.scala 102:19]
  wire  m_748_io_x2; // @[MUL.scala 102:19]
  wire  m_748_io_x3; // @[MUL.scala 102:19]
  wire  m_748_io_s; // @[MUL.scala 102:19]
  wire  m_748_io_cout; // @[MUL.scala 102:19]
  wire  m_749_io_x1; // @[MUL.scala 102:19]
  wire  m_749_io_x2; // @[MUL.scala 102:19]
  wire  m_749_io_x3; // @[MUL.scala 102:19]
  wire  m_749_io_s; // @[MUL.scala 102:19]
  wire  m_749_io_cout; // @[MUL.scala 102:19]
  wire  m_750_io_x1; // @[MUL.scala 102:19]
  wire  m_750_io_x2; // @[MUL.scala 102:19]
  wire  m_750_io_x3; // @[MUL.scala 102:19]
  wire  m_750_io_s; // @[MUL.scala 102:19]
  wire  m_750_io_cout; // @[MUL.scala 102:19]
  wire  m_751_io_x1; // @[MUL.scala 102:19]
  wire  m_751_io_x2; // @[MUL.scala 102:19]
  wire  m_751_io_x3; // @[MUL.scala 102:19]
  wire  m_751_io_s; // @[MUL.scala 102:19]
  wire  m_751_io_cout; // @[MUL.scala 102:19]
  wire  m_752_io_x1; // @[MUL.scala 102:19]
  wire  m_752_io_x2; // @[MUL.scala 102:19]
  wire  m_752_io_x3; // @[MUL.scala 102:19]
  wire  m_752_io_s; // @[MUL.scala 102:19]
  wire  m_752_io_cout; // @[MUL.scala 102:19]
  wire  m_753_io_x1; // @[MUL.scala 102:19]
  wire  m_753_io_x2; // @[MUL.scala 102:19]
  wire  m_753_io_x3; // @[MUL.scala 102:19]
  wire  m_753_io_s; // @[MUL.scala 102:19]
  wire  m_753_io_cout; // @[MUL.scala 102:19]
  wire  m_754_io_x1; // @[MUL.scala 102:19]
  wire  m_754_io_x2; // @[MUL.scala 102:19]
  wire  m_754_io_x3; // @[MUL.scala 102:19]
  wire  m_754_io_s; // @[MUL.scala 102:19]
  wire  m_754_io_cout; // @[MUL.scala 102:19]
  wire  m_755_io_x1; // @[MUL.scala 102:19]
  wire  m_755_io_x2; // @[MUL.scala 102:19]
  wire  m_755_io_x3; // @[MUL.scala 102:19]
  wire  m_755_io_s; // @[MUL.scala 102:19]
  wire  m_755_io_cout; // @[MUL.scala 102:19]
  wire  m_756_io_x1; // @[MUL.scala 102:19]
  wire  m_756_io_x2; // @[MUL.scala 102:19]
  wire  m_756_io_x3; // @[MUL.scala 102:19]
  wire  m_756_io_s; // @[MUL.scala 102:19]
  wire  m_756_io_cout; // @[MUL.scala 102:19]
  wire  m_757_io_x1; // @[MUL.scala 102:19]
  wire  m_757_io_x2; // @[MUL.scala 102:19]
  wire  m_757_io_x3; // @[MUL.scala 102:19]
  wire  m_757_io_s; // @[MUL.scala 102:19]
  wire  m_757_io_cout; // @[MUL.scala 102:19]
  wire  m_758_io_x1; // @[MUL.scala 102:19]
  wire  m_758_io_x2; // @[MUL.scala 102:19]
  wire  m_758_io_x3; // @[MUL.scala 102:19]
  wire  m_758_io_s; // @[MUL.scala 102:19]
  wire  m_758_io_cout; // @[MUL.scala 102:19]
  wire  m_759_io_x1; // @[MUL.scala 102:19]
  wire  m_759_io_x2; // @[MUL.scala 102:19]
  wire  m_759_io_x3; // @[MUL.scala 102:19]
  wire  m_759_io_s; // @[MUL.scala 102:19]
  wire  m_759_io_cout; // @[MUL.scala 102:19]
  wire  m_760_io_x1; // @[MUL.scala 102:19]
  wire  m_760_io_x2; // @[MUL.scala 102:19]
  wire  m_760_io_x3; // @[MUL.scala 102:19]
  wire  m_760_io_s; // @[MUL.scala 102:19]
  wire  m_760_io_cout; // @[MUL.scala 102:19]
  wire  m_761_io_x1; // @[MUL.scala 102:19]
  wire  m_761_io_x2; // @[MUL.scala 102:19]
  wire  m_761_io_x3; // @[MUL.scala 102:19]
  wire  m_761_io_s; // @[MUL.scala 102:19]
  wire  m_761_io_cout; // @[MUL.scala 102:19]
  wire  m_762_io_in_0; // @[MUL.scala 124:19]
  wire  m_762_io_in_1; // @[MUL.scala 124:19]
  wire  m_762_io_out_0; // @[MUL.scala 124:19]
  wire  m_762_io_out_1; // @[MUL.scala 124:19]
  wire  m_763_io_x1; // @[MUL.scala 102:19]
  wire  m_763_io_x2; // @[MUL.scala 102:19]
  wire  m_763_io_x3; // @[MUL.scala 102:19]
  wire  m_763_io_s; // @[MUL.scala 102:19]
  wire  m_763_io_cout; // @[MUL.scala 102:19]
  wire  m_764_io_x1; // @[MUL.scala 102:19]
  wire  m_764_io_x2; // @[MUL.scala 102:19]
  wire  m_764_io_x3; // @[MUL.scala 102:19]
  wire  m_764_io_s; // @[MUL.scala 102:19]
  wire  m_764_io_cout; // @[MUL.scala 102:19]
  wire  m_765_io_x1; // @[MUL.scala 102:19]
  wire  m_765_io_x2; // @[MUL.scala 102:19]
  wire  m_765_io_x3; // @[MUL.scala 102:19]
  wire  m_765_io_s; // @[MUL.scala 102:19]
  wire  m_765_io_cout; // @[MUL.scala 102:19]
  wire  m_766_io_in_0; // @[MUL.scala 124:19]
  wire  m_766_io_in_1; // @[MUL.scala 124:19]
  wire  m_766_io_out_0; // @[MUL.scala 124:19]
  wire  m_766_io_out_1; // @[MUL.scala 124:19]
  wire  m_767_io_x1; // @[MUL.scala 102:19]
  wire  m_767_io_x2; // @[MUL.scala 102:19]
  wire  m_767_io_x3; // @[MUL.scala 102:19]
  wire  m_767_io_s; // @[MUL.scala 102:19]
  wire  m_767_io_cout; // @[MUL.scala 102:19]
  wire  m_768_io_x1; // @[MUL.scala 102:19]
  wire  m_768_io_x2; // @[MUL.scala 102:19]
  wire  m_768_io_x3; // @[MUL.scala 102:19]
  wire  m_768_io_s; // @[MUL.scala 102:19]
  wire  m_768_io_cout; // @[MUL.scala 102:19]
  wire  m_769_io_x1; // @[MUL.scala 102:19]
  wire  m_769_io_x2; // @[MUL.scala 102:19]
  wire  m_769_io_x3; // @[MUL.scala 102:19]
  wire  m_769_io_s; // @[MUL.scala 102:19]
  wire  m_769_io_cout; // @[MUL.scala 102:19]
  wire  m_770_io_x1; // @[MUL.scala 102:19]
  wire  m_770_io_x2; // @[MUL.scala 102:19]
  wire  m_770_io_x3; // @[MUL.scala 102:19]
  wire  m_770_io_s; // @[MUL.scala 102:19]
  wire  m_770_io_cout; // @[MUL.scala 102:19]
  wire  m_771_io_x1; // @[MUL.scala 102:19]
  wire  m_771_io_x2; // @[MUL.scala 102:19]
  wire  m_771_io_x3; // @[MUL.scala 102:19]
  wire  m_771_io_s; // @[MUL.scala 102:19]
  wire  m_771_io_cout; // @[MUL.scala 102:19]
  wire  m_772_io_x1; // @[MUL.scala 102:19]
  wire  m_772_io_x2; // @[MUL.scala 102:19]
  wire  m_772_io_x3; // @[MUL.scala 102:19]
  wire  m_772_io_s; // @[MUL.scala 102:19]
  wire  m_772_io_cout; // @[MUL.scala 102:19]
  wire  m_773_io_x1; // @[MUL.scala 102:19]
  wire  m_773_io_x2; // @[MUL.scala 102:19]
  wire  m_773_io_x3; // @[MUL.scala 102:19]
  wire  m_773_io_s; // @[MUL.scala 102:19]
  wire  m_773_io_cout; // @[MUL.scala 102:19]
  wire  m_774_io_x1; // @[MUL.scala 102:19]
  wire  m_774_io_x2; // @[MUL.scala 102:19]
  wire  m_774_io_x3; // @[MUL.scala 102:19]
  wire  m_774_io_s; // @[MUL.scala 102:19]
  wire  m_774_io_cout; // @[MUL.scala 102:19]
  wire  m_775_io_x1; // @[MUL.scala 102:19]
  wire  m_775_io_x2; // @[MUL.scala 102:19]
  wire  m_775_io_x3; // @[MUL.scala 102:19]
  wire  m_775_io_s; // @[MUL.scala 102:19]
  wire  m_775_io_cout; // @[MUL.scala 102:19]
  wire  m_776_io_x1; // @[MUL.scala 102:19]
  wire  m_776_io_x2; // @[MUL.scala 102:19]
  wire  m_776_io_x3; // @[MUL.scala 102:19]
  wire  m_776_io_s; // @[MUL.scala 102:19]
  wire  m_776_io_cout; // @[MUL.scala 102:19]
  wire  m_777_io_x1; // @[MUL.scala 102:19]
  wire  m_777_io_x2; // @[MUL.scala 102:19]
  wire  m_777_io_x3; // @[MUL.scala 102:19]
  wire  m_777_io_s; // @[MUL.scala 102:19]
  wire  m_777_io_cout; // @[MUL.scala 102:19]
  wire  m_778_io_x1; // @[MUL.scala 102:19]
  wire  m_778_io_x2; // @[MUL.scala 102:19]
  wire  m_778_io_x3; // @[MUL.scala 102:19]
  wire  m_778_io_s; // @[MUL.scala 102:19]
  wire  m_778_io_cout; // @[MUL.scala 102:19]
  wire  m_779_io_x1; // @[MUL.scala 102:19]
  wire  m_779_io_x2; // @[MUL.scala 102:19]
  wire  m_779_io_x3; // @[MUL.scala 102:19]
  wire  m_779_io_s; // @[MUL.scala 102:19]
  wire  m_779_io_cout; // @[MUL.scala 102:19]
  wire  m_780_io_x1; // @[MUL.scala 102:19]
  wire  m_780_io_x2; // @[MUL.scala 102:19]
  wire  m_780_io_x3; // @[MUL.scala 102:19]
  wire  m_780_io_s; // @[MUL.scala 102:19]
  wire  m_780_io_cout; // @[MUL.scala 102:19]
  wire  m_781_io_in_0; // @[MUL.scala 124:19]
  wire  m_781_io_in_1; // @[MUL.scala 124:19]
  wire  m_781_io_out_0; // @[MUL.scala 124:19]
  wire  m_781_io_out_1; // @[MUL.scala 124:19]
  wire  m_782_io_x1; // @[MUL.scala 102:19]
  wire  m_782_io_x2; // @[MUL.scala 102:19]
  wire  m_782_io_x3; // @[MUL.scala 102:19]
  wire  m_782_io_s; // @[MUL.scala 102:19]
  wire  m_782_io_cout; // @[MUL.scala 102:19]
  wire  m_783_io_x1; // @[MUL.scala 102:19]
  wire  m_783_io_x2; // @[MUL.scala 102:19]
  wire  m_783_io_x3; // @[MUL.scala 102:19]
  wire  m_783_io_s; // @[MUL.scala 102:19]
  wire  m_783_io_cout; // @[MUL.scala 102:19]
  wire  m_784_io_in_0; // @[MUL.scala 124:19]
  wire  m_784_io_in_1; // @[MUL.scala 124:19]
  wire  m_784_io_out_0; // @[MUL.scala 124:19]
  wire  m_784_io_out_1; // @[MUL.scala 124:19]
  wire  m_785_io_x1; // @[MUL.scala 102:19]
  wire  m_785_io_x2; // @[MUL.scala 102:19]
  wire  m_785_io_x3; // @[MUL.scala 102:19]
  wire  m_785_io_s; // @[MUL.scala 102:19]
  wire  m_785_io_cout; // @[MUL.scala 102:19]
  wire  m_786_io_x1; // @[MUL.scala 102:19]
  wire  m_786_io_x2; // @[MUL.scala 102:19]
  wire  m_786_io_x3; // @[MUL.scala 102:19]
  wire  m_786_io_s; // @[MUL.scala 102:19]
  wire  m_786_io_cout; // @[MUL.scala 102:19]
  wire  m_787_io_x1; // @[MUL.scala 102:19]
  wire  m_787_io_x2; // @[MUL.scala 102:19]
  wire  m_787_io_x3; // @[MUL.scala 102:19]
  wire  m_787_io_s; // @[MUL.scala 102:19]
  wire  m_787_io_cout; // @[MUL.scala 102:19]
  wire  m_788_io_x1; // @[MUL.scala 102:19]
  wire  m_788_io_x2; // @[MUL.scala 102:19]
  wire  m_788_io_x3; // @[MUL.scala 102:19]
  wire  m_788_io_s; // @[MUL.scala 102:19]
  wire  m_788_io_cout; // @[MUL.scala 102:19]
  wire  m_789_io_x1; // @[MUL.scala 102:19]
  wire  m_789_io_x2; // @[MUL.scala 102:19]
  wire  m_789_io_x3; // @[MUL.scala 102:19]
  wire  m_789_io_s; // @[MUL.scala 102:19]
  wire  m_789_io_cout; // @[MUL.scala 102:19]
  wire  m_790_io_x1; // @[MUL.scala 102:19]
  wire  m_790_io_x2; // @[MUL.scala 102:19]
  wire  m_790_io_x3; // @[MUL.scala 102:19]
  wire  m_790_io_s; // @[MUL.scala 102:19]
  wire  m_790_io_cout; // @[MUL.scala 102:19]
  wire  m_791_io_x1; // @[MUL.scala 102:19]
  wire  m_791_io_x2; // @[MUL.scala 102:19]
  wire  m_791_io_x3; // @[MUL.scala 102:19]
  wire  m_791_io_s; // @[MUL.scala 102:19]
  wire  m_791_io_cout; // @[MUL.scala 102:19]
  wire  m_792_io_x1; // @[MUL.scala 102:19]
  wire  m_792_io_x2; // @[MUL.scala 102:19]
  wire  m_792_io_x3; // @[MUL.scala 102:19]
  wire  m_792_io_s; // @[MUL.scala 102:19]
  wire  m_792_io_cout; // @[MUL.scala 102:19]
  wire  m_793_io_x1; // @[MUL.scala 102:19]
  wire  m_793_io_x2; // @[MUL.scala 102:19]
  wire  m_793_io_x3; // @[MUL.scala 102:19]
  wire  m_793_io_s; // @[MUL.scala 102:19]
  wire  m_793_io_cout; // @[MUL.scala 102:19]
  wire  m_794_io_in_0; // @[MUL.scala 124:19]
  wire  m_794_io_in_1; // @[MUL.scala 124:19]
  wire  m_794_io_out_0; // @[MUL.scala 124:19]
  wire  m_794_io_out_1; // @[MUL.scala 124:19]
  wire  m_795_io_x1; // @[MUL.scala 102:19]
  wire  m_795_io_x2; // @[MUL.scala 102:19]
  wire  m_795_io_x3; // @[MUL.scala 102:19]
  wire  m_795_io_s; // @[MUL.scala 102:19]
  wire  m_795_io_cout; // @[MUL.scala 102:19]
  wire  m_796_io_in_0; // @[MUL.scala 124:19]
  wire  m_796_io_in_1; // @[MUL.scala 124:19]
  wire  m_796_io_out_0; // @[MUL.scala 124:19]
  wire  m_796_io_out_1; // @[MUL.scala 124:19]
  wire  m_797_io_x1; // @[MUL.scala 102:19]
  wire  m_797_io_x2; // @[MUL.scala 102:19]
  wire  m_797_io_x3; // @[MUL.scala 102:19]
  wire  m_797_io_s; // @[MUL.scala 102:19]
  wire  m_797_io_cout; // @[MUL.scala 102:19]
  wire  m_798_io_x1; // @[MUL.scala 102:19]
  wire  m_798_io_x2; // @[MUL.scala 102:19]
  wire  m_798_io_x3; // @[MUL.scala 102:19]
  wire  m_798_io_s; // @[MUL.scala 102:19]
  wire  m_798_io_cout; // @[MUL.scala 102:19]
  wire  m_799_io_x1; // @[MUL.scala 102:19]
  wire  m_799_io_x2; // @[MUL.scala 102:19]
  wire  m_799_io_x3; // @[MUL.scala 102:19]
  wire  m_799_io_s; // @[MUL.scala 102:19]
  wire  m_799_io_cout; // @[MUL.scala 102:19]
  wire  m_800_io_x1; // @[MUL.scala 102:19]
  wire  m_800_io_x2; // @[MUL.scala 102:19]
  wire  m_800_io_x3; // @[MUL.scala 102:19]
  wire  m_800_io_s; // @[MUL.scala 102:19]
  wire  m_800_io_cout; // @[MUL.scala 102:19]
  wire  m_801_io_in_0; // @[MUL.scala 124:19]
  wire  m_801_io_in_1; // @[MUL.scala 124:19]
  wire  m_801_io_out_0; // @[MUL.scala 124:19]
  wire  m_801_io_out_1; // @[MUL.scala 124:19]
  wire  m_802_io_in_0; // @[MUL.scala 124:19]
  wire  m_802_io_in_1; // @[MUL.scala 124:19]
  wire  m_802_io_out_0; // @[MUL.scala 124:19]
  wire  m_802_io_out_1; // @[MUL.scala 124:19]
  wire  m_803_io_in_0; // @[MUL.scala 124:19]
  wire  m_803_io_in_1; // @[MUL.scala 124:19]
  wire  m_803_io_out_0; // @[MUL.scala 124:19]
  wire  m_803_io_out_1; // @[MUL.scala 124:19]
  wire  m_804_io_in_0; // @[MUL.scala 124:19]
  wire  m_804_io_in_1; // @[MUL.scala 124:19]
  wire  m_804_io_out_0; // @[MUL.scala 124:19]
  wire  m_804_io_out_1; // @[MUL.scala 124:19]
  wire  m_805_io_in_0; // @[MUL.scala 124:19]
  wire  m_805_io_in_1; // @[MUL.scala 124:19]
  wire  m_805_io_out_0; // @[MUL.scala 124:19]
  wire  m_805_io_out_1; // @[MUL.scala 124:19]
  wire  m_806_io_x1; // @[MUL.scala 102:19]
  wire  m_806_io_x2; // @[MUL.scala 102:19]
  wire  m_806_io_x3; // @[MUL.scala 102:19]
  wire  m_806_io_s; // @[MUL.scala 102:19]
  wire  m_806_io_cout; // @[MUL.scala 102:19]
  wire  m_807_io_x1; // @[MUL.scala 102:19]
  wire  m_807_io_x2; // @[MUL.scala 102:19]
  wire  m_807_io_x3; // @[MUL.scala 102:19]
  wire  m_807_io_s; // @[MUL.scala 102:19]
  wire  m_807_io_cout; // @[MUL.scala 102:19]
  wire  m_808_io_x1; // @[MUL.scala 102:19]
  wire  m_808_io_x2; // @[MUL.scala 102:19]
  wire  m_808_io_x3; // @[MUL.scala 102:19]
  wire  m_808_io_s; // @[MUL.scala 102:19]
  wire  m_808_io_cout; // @[MUL.scala 102:19]
  wire  m_809_io_x1; // @[MUL.scala 102:19]
  wire  m_809_io_x2; // @[MUL.scala 102:19]
  wire  m_809_io_x3; // @[MUL.scala 102:19]
  wire  m_809_io_s; // @[MUL.scala 102:19]
  wire  m_809_io_cout; // @[MUL.scala 102:19]
  wire  m_810_io_x1; // @[MUL.scala 102:19]
  wire  m_810_io_x2; // @[MUL.scala 102:19]
  wire  m_810_io_x3; // @[MUL.scala 102:19]
  wire  m_810_io_s; // @[MUL.scala 102:19]
  wire  m_810_io_cout; // @[MUL.scala 102:19]
  wire  m_811_io_x1; // @[MUL.scala 102:19]
  wire  m_811_io_x2; // @[MUL.scala 102:19]
  wire  m_811_io_x3; // @[MUL.scala 102:19]
  wire  m_811_io_s; // @[MUL.scala 102:19]
  wire  m_811_io_cout; // @[MUL.scala 102:19]
  wire  m_812_io_x1; // @[MUL.scala 102:19]
  wire  m_812_io_x2; // @[MUL.scala 102:19]
  wire  m_812_io_x3; // @[MUL.scala 102:19]
  wire  m_812_io_s; // @[MUL.scala 102:19]
  wire  m_812_io_cout; // @[MUL.scala 102:19]
  wire  m_813_io_in_0; // @[MUL.scala 124:19]
  wire  m_813_io_in_1; // @[MUL.scala 124:19]
  wire  m_813_io_out_0; // @[MUL.scala 124:19]
  wire  m_813_io_out_1; // @[MUL.scala 124:19]
  wire  m_814_io_x1; // @[MUL.scala 102:19]
  wire  m_814_io_x2; // @[MUL.scala 102:19]
  wire  m_814_io_x3; // @[MUL.scala 102:19]
  wire  m_814_io_s; // @[MUL.scala 102:19]
  wire  m_814_io_cout; // @[MUL.scala 102:19]
  wire  m_815_io_in_0; // @[MUL.scala 124:19]
  wire  m_815_io_in_1; // @[MUL.scala 124:19]
  wire  m_815_io_out_0; // @[MUL.scala 124:19]
  wire  m_815_io_out_1; // @[MUL.scala 124:19]
  wire  m_816_io_x1; // @[MUL.scala 102:19]
  wire  m_816_io_x2; // @[MUL.scala 102:19]
  wire  m_816_io_x3; // @[MUL.scala 102:19]
  wire  m_816_io_s; // @[MUL.scala 102:19]
  wire  m_816_io_cout; // @[MUL.scala 102:19]
  wire  m_817_io_in_0; // @[MUL.scala 124:19]
  wire  m_817_io_in_1; // @[MUL.scala 124:19]
  wire  m_817_io_out_0; // @[MUL.scala 124:19]
  wire  m_817_io_out_1; // @[MUL.scala 124:19]
  wire  m_818_io_x1; // @[MUL.scala 102:19]
  wire  m_818_io_x2; // @[MUL.scala 102:19]
  wire  m_818_io_x3; // @[MUL.scala 102:19]
  wire  m_818_io_s; // @[MUL.scala 102:19]
  wire  m_818_io_cout; // @[MUL.scala 102:19]
  wire  m_819_io_x1; // @[MUL.scala 102:19]
  wire  m_819_io_x2; // @[MUL.scala 102:19]
  wire  m_819_io_x3; // @[MUL.scala 102:19]
  wire  m_819_io_s; // @[MUL.scala 102:19]
  wire  m_819_io_cout; // @[MUL.scala 102:19]
  wire  m_820_io_x1; // @[MUL.scala 102:19]
  wire  m_820_io_x2; // @[MUL.scala 102:19]
  wire  m_820_io_x3; // @[MUL.scala 102:19]
  wire  m_820_io_s; // @[MUL.scala 102:19]
  wire  m_820_io_cout; // @[MUL.scala 102:19]
  wire  m_821_io_x1; // @[MUL.scala 102:19]
  wire  m_821_io_x2; // @[MUL.scala 102:19]
  wire  m_821_io_x3; // @[MUL.scala 102:19]
  wire  m_821_io_s; // @[MUL.scala 102:19]
  wire  m_821_io_cout; // @[MUL.scala 102:19]
  wire  m_822_io_x1; // @[MUL.scala 102:19]
  wire  m_822_io_x2; // @[MUL.scala 102:19]
  wire  m_822_io_x3; // @[MUL.scala 102:19]
  wire  m_822_io_s; // @[MUL.scala 102:19]
  wire  m_822_io_cout; // @[MUL.scala 102:19]
  wire  m_823_io_x1; // @[MUL.scala 102:19]
  wire  m_823_io_x2; // @[MUL.scala 102:19]
  wire  m_823_io_x3; // @[MUL.scala 102:19]
  wire  m_823_io_s; // @[MUL.scala 102:19]
  wire  m_823_io_cout; // @[MUL.scala 102:19]
  wire  m_824_io_x1; // @[MUL.scala 102:19]
  wire  m_824_io_x2; // @[MUL.scala 102:19]
  wire  m_824_io_x3; // @[MUL.scala 102:19]
  wire  m_824_io_s; // @[MUL.scala 102:19]
  wire  m_824_io_cout; // @[MUL.scala 102:19]
  wire  m_825_io_x1; // @[MUL.scala 102:19]
  wire  m_825_io_x2; // @[MUL.scala 102:19]
  wire  m_825_io_x3; // @[MUL.scala 102:19]
  wire  m_825_io_s; // @[MUL.scala 102:19]
  wire  m_825_io_cout; // @[MUL.scala 102:19]
  wire  m_826_io_x1; // @[MUL.scala 102:19]
  wire  m_826_io_x2; // @[MUL.scala 102:19]
  wire  m_826_io_x3; // @[MUL.scala 102:19]
  wire  m_826_io_s; // @[MUL.scala 102:19]
  wire  m_826_io_cout; // @[MUL.scala 102:19]
  wire  m_827_io_x1; // @[MUL.scala 102:19]
  wire  m_827_io_x2; // @[MUL.scala 102:19]
  wire  m_827_io_x3; // @[MUL.scala 102:19]
  wire  m_827_io_s; // @[MUL.scala 102:19]
  wire  m_827_io_cout; // @[MUL.scala 102:19]
  wire  m_828_io_x1; // @[MUL.scala 102:19]
  wire  m_828_io_x2; // @[MUL.scala 102:19]
  wire  m_828_io_x3; // @[MUL.scala 102:19]
  wire  m_828_io_s; // @[MUL.scala 102:19]
  wire  m_828_io_cout; // @[MUL.scala 102:19]
  wire  m_829_io_x1; // @[MUL.scala 102:19]
  wire  m_829_io_x2; // @[MUL.scala 102:19]
  wire  m_829_io_x3; // @[MUL.scala 102:19]
  wire  m_829_io_s; // @[MUL.scala 102:19]
  wire  m_829_io_cout; // @[MUL.scala 102:19]
  wire  m_830_io_x1; // @[MUL.scala 102:19]
  wire  m_830_io_x2; // @[MUL.scala 102:19]
  wire  m_830_io_x3; // @[MUL.scala 102:19]
  wire  m_830_io_s; // @[MUL.scala 102:19]
  wire  m_830_io_cout; // @[MUL.scala 102:19]
  wire  m_831_io_x1; // @[MUL.scala 102:19]
  wire  m_831_io_x2; // @[MUL.scala 102:19]
  wire  m_831_io_x3; // @[MUL.scala 102:19]
  wire  m_831_io_s; // @[MUL.scala 102:19]
  wire  m_831_io_cout; // @[MUL.scala 102:19]
  wire  m_832_io_in_0; // @[MUL.scala 124:19]
  wire  m_832_io_in_1; // @[MUL.scala 124:19]
  wire  m_832_io_out_0; // @[MUL.scala 124:19]
  wire  m_832_io_out_1; // @[MUL.scala 124:19]
  wire  m_833_io_x1; // @[MUL.scala 102:19]
  wire  m_833_io_x2; // @[MUL.scala 102:19]
  wire  m_833_io_x3; // @[MUL.scala 102:19]
  wire  m_833_io_s; // @[MUL.scala 102:19]
  wire  m_833_io_cout; // @[MUL.scala 102:19]
  wire  m_834_io_x1; // @[MUL.scala 102:19]
  wire  m_834_io_x2; // @[MUL.scala 102:19]
  wire  m_834_io_x3; // @[MUL.scala 102:19]
  wire  m_834_io_s; // @[MUL.scala 102:19]
  wire  m_834_io_cout; // @[MUL.scala 102:19]
  wire  m_835_io_in_0; // @[MUL.scala 124:19]
  wire  m_835_io_in_1; // @[MUL.scala 124:19]
  wire  m_835_io_out_0; // @[MUL.scala 124:19]
  wire  m_835_io_out_1; // @[MUL.scala 124:19]
  wire  m_836_io_x1; // @[MUL.scala 102:19]
  wire  m_836_io_x2; // @[MUL.scala 102:19]
  wire  m_836_io_x3; // @[MUL.scala 102:19]
  wire  m_836_io_s; // @[MUL.scala 102:19]
  wire  m_836_io_cout; // @[MUL.scala 102:19]
  wire  m_837_io_x1; // @[MUL.scala 102:19]
  wire  m_837_io_x2; // @[MUL.scala 102:19]
  wire  m_837_io_x3; // @[MUL.scala 102:19]
  wire  m_837_io_s; // @[MUL.scala 102:19]
  wire  m_837_io_cout; // @[MUL.scala 102:19]
  wire  m_838_io_in_0; // @[MUL.scala 124:19]
  wire  m_838_io_in_1; // @[MUL.scala 124:19]
  wire  m_838_io_out_0; // @[MUL.scala 124:19]
  wire  m_838_io_out_1; // @[MUL.scala 124:19]
  wire  m_839_io_x1; // @[MUL.scala 102:19]
  wire  m_839_io_x2; // @[MUL.scala 102:19]
  wire  m_839_io_x3; // @[MUL.scala 102:19]
  wire  m_839_io_s; // @[MUL.scala 102:19]
  wire  m_839_io_cout; // @[MUL.scala 102:19]
  wire  m_840_io_x1; // @[MUL.scala 102:19]
  wire  m_840_io_x2; // @[MUL.scala 102:19]
  wire  m_840_io_x3; // @[MUL.scala 102:19]
  wire  m_840_io_s; // @[MUL.scala 102:19]
  wire  m_840_io_cout; // @[MUL.scala 102:19]
  wire  m_841_io_x1; // @[MUL.scala 102:19]
  wire  m_841_io_x2; // @[MUL.scala 102:19]
  wire  m_841_io_x3; // @[MUL.scala 102:19]
  wire  m_841_io_s; // @[MUL.scala 102:19]
  wire  m_841_io_cout; // @[MUL.scala 102:19]
  wire  m_842_io_x1; // @[MUL.scala 102:19]
  wire  m_842_io_x2; // @[MUL.scala 102:19]
  wire  m_842_io_x3; // @[MUL.scala 102:19]
  wire  m_842_io_s; // @[MUL.scala 102:19]
  wire  m_842_io_cout; // @[MUL.scala 102:19]
  wire  m_843_io_x1; // @[MUL.scala 102:19]
  wire  m_843_io_x2; // @[MUL.scala 102:19]
  wire  m_843_io_x3; // @[MUL.scala 102:19]
  wire  m_843_io_s; // @[MUL.scala 102:19]
  wire  m_843_io_cout; // @[MUL.scala 102:19]
  wire  m_844_io_x1; // @[MUL.scala 102:19]
  wire  m_844_io_x2; // @[MUL.scala 102:19]
  wire  m_844_io_x3; // @[MUL.scala 102:19]
  wire  m_844_io_s; // @[MUL.scala 102:19]
  wire  m_844_io_cout; // @[MUL.scala 102:19]
  wire  m_845_io_x1; // @[MUL.scala 102:19]
  wire  m_845_io_x2; // @[MUL.scala 102:19]
  wire  m_845_io_x3; // @[MUL.scala 102:19]
  wire  m_845_io_s; // @[MUL.scala 102:19]
  wire  m_845_io_cout; // @[MUL.scala 102:19]
  wire  m_846_io_x1; // @[MUL.scala 102:19]
  wire  m_846_io_x2; // @[MUL.scala 102:19]
  wire  m_846_io_x3; // @[MUL.scala 102:19]
  wire  m_846_io_s; // @[MUL.scala 102:19]
  wire  m_846_io_cout; // @[MUL.scala 102:19]
  wire  m_847_io_x1; // @[MUL.scala 102:19]
  wire  m_847_io_x2; // @[MUL.scala 102:19]
  wire  m_847_io_x3; // @[MUL.scala 102:19]
  wire  m_847_io_s; // @[MUL.scala 102:19]
  wire  m_847_io_cout; // @[MUL.scala 102:19]
  wire  m_848_io_x1; // @[MUL.scala 102:19]
  wire  m_848_io_x2; // @[MUL.scala 102:19]
  wire  m_848_io_x3; // @[MUL.scala 102:19]
  wire  m_848_io_s; // @[MUL.scala 102:19]
  wire  m_848_io_cout; // @[MUL.scala 102:19]
  wire  m_849_io_x1; // @[MUL.scala 102:19]
  wire  m_849_io_x2; // @[MUL.scala 102:19]
  wire  m_849_io_x3; // @[MUL.scala 102:19]
  wire  m_849_io_s; // @[MUL.scala 102:19]
  wire  m_849_io_cout; // @[MUL.scala 102:19]
  wire  m_850_io_x1; // @[MUL.scala 102:19]
  wire  m_850_io_x2; // @[MUL.scala 102:19]
  wire  m_850_io_x3; // @[MUL.scala 102:19]
  wire  m_850_io_s; // @[MUL.scala 102:19]
  wire  m_850_io_cout; // @[MUL.scala 102:19]
  wire  m_851_io_x1; // @[MUL.scala 102:19]
  wire  m_851_io_x2; // @[MUL.scala 102:19]
  wire  m_851_io_x3; // @[MUL.scala 102:19]
  wire  m_851_io_s; // @[MUL.scala 102:19]
  wire  m_851_io_cout; // @[MUL.scala 102:19]
  wire  m_852_io_x1; // @[MUL.scala 102:19]
  wire  m_852_io_x2; // @[MUL.scala 102:19]
  wire  m_852_io_x3; // @[MUL.scala 102:19]
  wire  m_852_io_s; // @[MUL.scala 102:19]
  wire  m_852_io_cout; // @[MUL.scala 102:19]
  wire  m_853_io_x1; // @[MUL.scala 102:19]
  wire  m_853_io_x2; // @[MUL.scala 102:19]
  wire  m_853_io_x3; // @[MUL.scala 102:19]
  wire  m_853_io_s; // @[MUL.scala 102:19]
  wire  m_853_io_cout; // @[MUL.scala 102:19]
  wire  m_854_io_x1; // @[MUL.scala 102:19]
  wire  m_854_io_x2; // @[MUL.scala 102:19]
  wire  m_854_io_x3; // @[MUL.scala 102:19]
  wire  m_854_io_s; // @[MUL.scala 102:19]
  wire  m_854_io_cout; // @[MUL.scala 102:19]
  wire  m_855_io_x1; // @[MUL.scala 102:19]
  wire  m_855_io_x2; // @[MUL.scala 102:19]
  wire  m_855_io_x3; // @[MUL.scala 102:19]
  wire  m_855_io_s; // @[MUL.scala 102:19]
  wire  m_855_io_cout; // @[MUL.scala 102:19]
  wire  m_856_io_x1; // @[MUL.scala 102:19]
  wire  m_856_io_x2; // @[MUL.scala 102:19]
  wire  m_856_io_x3; // @[MUL.scala 102:19]
  wire  m_856_io_s; // @[MUL.scala 102:19]
  wire  m_856_io_cout; // @[MUL.scala 102:19]
  wire  m_857_io_x1; // @[MUL.scala 102:19]
  wire  m_857_io_x2; // @[MUL.scala 102:19]
  wire  m_857_io_x3; // @[MUL.scala 102:19]
  wire  m_857_io_s; // @[MUL.scala 102:19]
  wire  m_857_io_cout; // @[MUL.scala 102:19]
  wire  m_858_io_x1; // @[MUL.scala 102:19]
  wire  m_858_io_x2; // @[MUL.scala 102:19]
  wire  m_858_io_x3; // @[MUL.scala 102:19]
  wire  m_858_io_s; // @[MUL.scala 102:19]
  wire  m_858_io_cout; // @[MUL.scala 102:19]
  wire  m_859_io_x1; // @[MUL.scala 102:19]
  wire  m_859_io_x2; // @[MUL.scala 102:19]
  wire  m_859_io_x3; // @[MUL.scala 102:19]
  wire  m_859_io_s; // @[MUL.scala 102:19]
  wire  m_859_io_cout; // @[MUL.scala 102:19]
  wire  m_860_io_in_0; // @[MUL.scala 124:19]
  wire  m_860_io_in_1; // @[MUL.scala 124:19]
  wire  m_860_io_out_0; // @[MUL.scala 124:19]
  wire  m_860_io_out_1; // @[MUL.scala 124:19]
  wire  m_861_io_x1; // @[MUL.scala 102:19]
  wire  m_861_io_x2; // @[MUL.scala 102:19]
  wire  m_861_io_x3; // @[MUL.scala 102:19]
  wire  m_861_io_s; // @[MUL.scala 102:19]
  wire  m_861_io_cout; // @[MUL.scala 102:19]
  wire  m_862_io_x1; // @[MUL.scala 102:19]
  wire  m_862_io_x2; // @[MUL.scala 102:19]
  wire  m_862_io_x3; // @[MUL.scala 102:19]
  wire  m_862_io_s; // @[MUL.scala 102:19]
  wire  m_862_io_cout; // @[MUL.scala 102:19]
  wire  m_863_io_x1; // @[MUL.scala 102:19]
  wire  m_863_io_x2; // @[MUL.scala 102:19]
  wire  m_863_io_x3; // @[MUL.scala 102:19]
  wire  m_863_io_s; // @[MUL.scala 102:19]
  wire  m_863_io_cout; // @[MUL.scala 102:19]
  wire  m_864_io_in_0; // @[MUL.scala 124:19]
  wire  m_864_io_in_1; // @[MUL.scala 124:19]
  wire  m_864_io_out_0; // @[MUL.scala 124:19]
  wire  m_864_io_out_1; // @[MUL.scala 124:19]
  wire  m_865_io_x1; // @[MUL.scala 102:19]
  wire  m_865_io_x2; // @[MUL.scala 102:19]
  wire  m_865_io_x3; // @[MUL.scala 102:19]
  wire  m_865_io_s; // @[MUL.scala 102:19]
  wire  m_865_io_cout; // @[MUL.scala 102:19]
  wire  m_866_io_x1; // @[MUL.scala 102:19]
  wire  m_866_io_x2; // @[MUL.scala 102:19]
  wire  m_866_io_x3; // @[MUL.scala 102:19]
  wire  m_866_io_s; // @[MUL.scala 102:19]
  wire  m_866_io_cout; // @[MUL.scala 102:19]
  wire  m_867_io_x1; // @[MUL.scala 102:19]
  wire  m_867_io_x2; // @[MUL.scala 102:19]
  wire  m_867_io_x3; // @[MUL.scala 102:19]
  wire  m_867_io_s; // @[MUL.scala 102:19]
  wire  m_867_io_cout; // @[MUL.scala 102:19]
  wire  m_868_io_in_0; // @[MUL.scala 124:19]
  wire  m_868_io_in_1; // @[MUL.scala 124:19]
  wire  m_868_io_out_0; // @[MUL.scala 124:19]
  wire  m_868_io_out_1; // @[MUL.scala 124:19]
  wire  m_869_io_x1; // @[MUL.scala 102:19]
  wire  m_869_io_x2; // @[MUL.scala 102:19]
  wire  m_869_io_x3; // @[MUL.scala 102:19]
  wire  m_869_io_s; // @[MUL.scala 102:19]
  wire  m_869_io_cout; // @[MUL.scala 102:19]
  wire  m_870_io_x1; // @[MUL.scala 102:19]
  wire  m_870_io_x2; // @[MUL.scala 102:19]
  wire  m_870_io_x3; // @[MUL.scala 102:19]
  wire  m_870_io_s; // @[MUL.scala 102:19]
  wire  m_870_io_cout; // @[MUL.scala 102:19]
  wire  m_871_io_x1; // @[MUL.scala 102:19]
  wire  m_871_io_x2; // @[MUL.scala 102:19]
  wire  m_871_io_x3; // @[MUL.scala 102:19]
  wire  m_871_io_s; // @[MUL.scala 102:19]
  wire  m_871_io_cout; // @[MUL.scala 102:19]
  wire  m_872_io_x1; // @[MUL.scala 102:19]
  wire  m_872_io_x2; // @[MUL.scala 102:19]
  wire  m_872_io_x3; // @[MUL.scala 102:19]
  wire  m_872_io_s; // @[MUL.scala 102:19]
  wire  m_872_io_cout; // @[MUL.scala 102:19]
  wire  m_873_io_x1; // @[MUL.scala 102:19]
  wire  m_873_io_x2; // @[MUL.scala 102:19]
  wire  m_873_io_x3; // @[MUL.scala 102:19]
  wire  m_873_io_s; // @[MUL.scala 102:19]
  wire  m_873_io_cout; // @[MUL.scala 102:19]
  wire  m_874_io_x1; // @[MUL.scala 102:19]
  wire  m_874_io_x2; // @[MUL.scala 102:19]
  wire  m_874_io_x3; // @[MUL.scala 102:19]
  wire  m_874_io_s; // @[MUL.scala 102:19]
  wire  m_874_io_cout; // @[MUL.scala 102:19]
  wire  m_875_io_x1; // @[MUL.scala 102:19]
  wire  m_875_io_x2; // @[MUL.scala 102:19]
  wire  m_875_io_x3; // @[MUL.scala 102:19]
  wire  m_875_io_s; // @[MUL.scala 102:19]
  wire  m_875_io_cout; // @[MUL.scala 102:19]
  wire  m_876_io_x1; // @[MUL.scala 102:19]
  wire  m_876_io_x2; // @[MUL.scala 102:19]
  wire  m_876_io_x3; // @[MUL.scala 102:19]
  wire  m_876_io_s; // @[MUL.scala 102:19]
  wire  m_876_io_cout; // @[MUL.scala 102:19]
  wire  m_877_io_x1; // @[MUL.scala 102:19]
  wire  m_877_io_x2; // @[MUL.scala 102:19]
  wire  m_877_io_x3; // @[MUL.scala 102:19]
  wire  m_877_io_s; // @[MUL.scala 102:19]
  wire  m_877_io_cout; // @[MUL.scala 102:19]
  wire  m_878_io_x1; // @[MUL.scala 102:19]
  wire  m_878_io_x2; // @[MUL.scala 102:19]
  wire  m_878_io_x3; // @[MUL.scala 102:19]
  wire  m_878_io_s; // @[MUL.scala 102:19]
  wire  m_878_io_cout; // @[MUL.scala 102:19]
  wire  m_879_io_x1; // @[MUL.scala 102:19]
  wire  m_879_io_x2; // @[MUL.scala 102:19]
  wire  m_879_io_x3; // @[MUL.scala 102:19]
  wire  m_879_io_s; // @[MUL.scala 102:19]
  wire  m_879_io_cout; // @[MUL.scala 102:19]
  wire  m_880_io_x1; // @[MUL.scala 102:19]
  wire  m_880_io_x2; // @[MUL.scala 102:19]
  wire  m_880_io_x3; // @[MUL.scala 102:19]
  wire  m_880_io_s; // @[MUL.scala 102:19]
  wire  m_880_io_cout; // @[MUL.scala 102:19]
  wire  m_881_io_x1; // @[MUL.scala 102:19]
  wire  m_881_io_x2; // @[MUL.scala 102:19]
  wire  m_881_io_x3; // @[MUL.scala 102:19]
  wire  m_881_io_s; // @[MUL.scala 102:19]
  wire  m_881_io_cout; // @[MUL.scala 102:19]
  wire  m_882_io_x1; // @[MUL.scala 102:19]
  wire  m_882_io_x2; // @[MUL.scala 102:19]
  wire  m_882_io_x3; // @[MUL.scala 102:19]
  wire  m_882_io_s; // @[MUL.scala 102:19]
  wire  m_882_io_cout; // @[MUL.scala 102:19]
  wire  m_883_io_x1; // @[MUL.scala 102:19]
  wire  m_883_io_x2; // @[MUL.scala 102:19]
  wire  m_883_io_x3; // @[MUL.scala 102:19]
  wire  m_883_io_s; // @[MUL.scala 102:19]
  wire  m_883_io_cout; // @[MUL.scala 102:19]
  wire  m_884_io_x1; // @[MUL.scala 102:19]
  wire  m_884_io_x2; // @[MUL.scala 102:19]
  wire  m_884_io_x3; // @[MUL.scala 102:19]
  wire  m_884_io_s; // @[MUL.scala 102:19]
  wire  m_884_io_cout; // @[MUL.scala 102:19]
  wire  m_885_io_x1; // @[MUL.scala 102:19]
  wire  m_885_io_x2; // @[MUL.scala 102:19]
  wire  m_885_io_x3; // @[MUL.scala 102:19]
  wire  m_885_io_s; // @[MUL.scala 102:19]
  wire  m_885_io_cout; // @[MUL.scala 102:19]
  wire  m_886_io_x1; // @[MUL.scala 102:19]
  wire  m_886_io_x2; // @[MUL.scala 102:19]
  wire  m_886_io_x3; // @[MUL.scala 102:19]
  wire  m_886_io_s; // @[MUL.scala 102:19]
  wire  m_886_io_cout; // @[MUL.scala 102:19]
  wire  m_887_io_x1; // @[MUL.scala 102:19]
  wire  m_887_io_x2; // @[MUL.scala 102:19]
  wire  m_887_io_x3; // @[MUL.scala 102:19]
  wire  m_887_io_s; // @[MUL.scala 102:19]
  wire  m_887_io_cout; // @[MUL.scala 102:19]
  wire  m_888_io_x1; // @[MUL.scala 102:19]
  wire  m_888_io_x2; // @[MUL.scala 102:19]
  wire  m_888_io_x3; // @[MUL.scala 102:19]
  wire  m_888_io_s; // @[MUL.scala 102:19]
  wire  m_888_io_cout; // @[MUL.scala 102:19]
  wire  m_889_io_x1; // @[MUL.scala 102:19]
  wire  m_889_io_x2; // @[MUL.scala 102:19]
  wire  m_889_io_x3; // @[MUL.scala 102:19]
  wire  m_889_io_s; // @[MUL.scala 102:19]
  wire  m_889_io_cout; // @[MUL.scala 102:19]
  wire  m_890_io_x1; // @[MUL.scala 102:19]
  wire  m_890_io_x2; // @[MUL.scala 102:19]
  wire  m_890_io_x3; // @[MUL.scala 102:19]
  wire  m_890_io_s; // @[MUL.scala 102:19]
  wire  m_890_io_cout; // @[MUL.scala 102:19]
  wire  m_891_io_x1; // @[MUL.scala 102:19]
  wire  m_891_io_x2; // @[MUL.scala 102:19]
  wire  m_891_io_x3; // @[MUL.scala 102:19]
  wire  m_891_io_s; // @[MUL.scala 102:19]
  wire  m_891_io_cout; // @[MUL.scala 102:19]
  wire  m_892_io_x1; // @[MUL.scala 102:19]
  wire  m_892_io_x2; // @[MUL.scala 102:19]
  wire  m_892_io_x3; // @[MUL.scala 102:19]
  wire  m_892_io_s; // @[MUL.scala 102:19]
  wire  m_892_io_cout; // @[MUL.scala 102:19]
  wire  m_893_io_x1; // @[MUL.scala 102:19]
  wire  m_893_io_x2; // @[MUL.scala 102:19]
  wire  m_893_io_x3; // @[MUL.scala 102:19]
  wire  m_893_io_s; // @[MUL.scala 102:19]
  wire  m_893_io_cout; // @[MUL.scala 102:19]
  wire  m_894_io_x1; // @[MUL.scala 102:19]
  wire  m_894_io_x2; // @[MUL.scala 102:19]
  wire  m_894_io_x3; // @[MUL.scala 102:19]
  wire  m_894_io_s; // @[MUL.scala 102:19]
  wire  m_894_io_cout; // @[MUL.scala 102:19]
  wire  m_895_io_x1; // @[MUL.scala 102:19]
  wire  m_895_io_x2; // @[MUL.scala 102:19]
  wire  m_895_io_x3; // @[MUL.scala 102:19]
  wire  m_895_io_s; // @[MUL.scala 102:19]
  wire  m_895_io_cout; // @[MUL.scala 102:19]
  wire  m_896_io_x1; // @[MUL.scala 102:19]
  wire  m_896_io_x2; // @[MUL.scala 102:19]
  wire  m_896_io_x3; // @[MUL.scala 102:19]
  wire  m_896_io_s; // @[MUL.scala 102:19]
  wire  m_896_io_cout; // @[MUL.scala 102:19]
  wire  m_897_io_in_0; // @[MUL.scala 124:19]
  wire  m_897_io_in_1; // @[MUL.scala 124:19]
  wire  m_897_io_out_0; // @[MUL.scala 124:19]
  wire  m_897_io_out_1; // @[MUL.scala 124:19]
  wire  m_898_io_x1; // @[MUL.scala 102:19]
  wire  m_898_io_x2; // @[MUL.scala 102:19]
  wire  m_898_io_x3; // @[MUL.scala 102:19]
  wire  m_898_io_s; // @[MUL.scala 102:19]
  wire  m_898_io_cout; // @[MUL.scala 102:19]
  wire  m_899_io_x1; // @[MUL.scala 102:19]
  wire  m_899_io_x2; // @[MUL.scala 102:19]
  wire  m_899_io_x3; // @[MUL.scala 102:19]
  wire  m_899_io_s; // @[MUL.scala 102:19]
  wire  m_899_io_cout; // @[MUL.scala 102:19]
  wire  m_900_io_x1; // @[MUL.scala 102:19]
  wire  m_900_io_x2; // @[MUL.scala 102:19]
  wire  m_900_io_x3; // @[MUL.scala 102:19]
  wire  m_900_io_s; // @[MUL.scala 102:19]
  wire  m_900_io_cout; // @[MUL.scala 102:19]
  wire  m_901_io_x1; // @[MUL.scala 102:19]
  wire  m_901_io_x2; // @[MUL.scala 102:19]
  wire  m_901_io_x3; // @[MUL.scala 102:19]
  wire  m_901_io_s; // @[MUL.scala 102:19]
  wire  m_901_io_cout; // @[MUL.scala 102:19]
  wire  m_902_io_in_0; // @[MUL.scala 124:19]
  wire  m_902_io_in_1; // @[MUL.scala 124:19]
  wire  m_902_io_out_0; // @[MUL.scala 124:19]
  wire  m_902_io_out_1; // @[MUL.scala 124:19]
  wire  m_903_io_x1; // @[MUL.scala 102:19]
  wire  m_903_io_x2; // @[MUL.scala 102:19]
  wire  m_903_io_x3; // @[MUL.scala 102:19]
  wire  m_903_io_s; // @[MUL.scala 102:19]
  wire  m_903_io_cout; // @[MUL.scala 102:19]
  wire  m_904_io_x1; // @[MUL.scala 102:19]
  wire  m_904_io_x2; // @[MUL.scala 102:19]
  wire  m_904_io_x3; // @[MUL.scala 102:19]
  wire  m_904_io_s; // @[MUL.scala 102:19]
  wire  m_904_io_cout; // @[MUL.scala 102:19]
  wire  m_905_io_x1; // @[MUL.scala 102:19]
  wire  m_905_io_x2; // @[MUL.scala 102:19]
  wire  m_905_io_x3; // @[MUL.scala 102:19]
  wire  m_905_io_s; // @[MUL.scala 102:19]
  wire  m_905_io_cout; // @[MUL.scala 102:19]
  wire  m_906_io_x1; // @[MUL.scala 102:19]
  wire  m_906_io_x2; // @[MUL.scala 102:19]
  wire  m_906_io_x3; // @[MUL.scala 102:19]
  wire  m_906_io_s; // @[MUL.scala 102:19]
  wire  m_906_io_cout; // @[MUL.scala 102:19]
  wire  m_907_io_in_0; // @[MUL.scala 124:19]
  wire  m_907_io_in_1; // @[MUL.scala 124:19]
  wire  m_907_io_out_0; // @[MUL.scala 124:19]
  wire  m_907_io_out_1; // @[MUL.scala 124:19]
  wire  m_908_io_x1; // @[MUL.scala 102:19]
  wire  m_908_io_x2; // @[MUL.scala 102:19]
  wire  m_908_io_x3; // @[MUL.scala 102:19]
  wire  m_908_io_s; // @[MUL.scala 102:19]
  wire  m_908_io_cout; // @[MUL.scala 102:19]
  wire  m_909_io_x1; // @[MUL.scala 102:19]
  wire  m_909_io_x2; // @[MUL.scala 102:19]
  wire  m_909_io_x3; // @[MUL.scala 102:19]
  wire  m_909_io_s; // @[MUL.scala 102:19]
  wire  m_909_io_cout; // @[MUL.scala 102:19]
  wire  m_910_io_x1; // @[MUL.scala 102:19]
  wire  m_910_io_x2; // @[MUL.scala 102:19]
  wire  m_910_io_x3; // @[MUL.scala 102:19]
  wire  m_910_io_s; // @[MUL.scala 102:19]
  wire  m_910_io_cout; // @[MUL.scala 102:19]
  wire  m_911_io_x1; // @[MUL.scala 102:19]
  wire  m_911_io_x2; // @[MUL.scala 102:19]
  wire  m_911_io_x3; // @[MUL.scala 102:19]
  wire  m_911_io_s; // @[MUL.scala 102:19]
  wire  m_911_io_cout; // @[MUL.scala 102:19]
  wire  m_912_io_x1; // @[MUL.scala 102:19]
  wire  m_912_io_x2; // @[MUL.scala 102:19]
  wire  m_912_io_x3; // @[MUL.scala 102:19]
  wire  m_912_io_s; // @[MUL.scala 102:19]
  wire  m_912_io_cout; // @[MUL.scala 102:19]
  wire  m_913_io_x1; // @[MUL.scala 102:19]
  wire  m_913_io_x2; // @[MUL.scala 102:19]
  wire  m_913_io_x3; // @[MUL.scala 102:19]
  wire  m_913_io_s; // @[MUL.scala 102:19]
  wire  m_913_io_cout; // @[MUL.scala 102:19]
  wire  m_914_io_x1; // @[MUL.scala 102:19]
  wire  m_914_io_x2; // @[MUL.scala 102:19]
  wire  m_914_io_x3; // @[MUL.scala 102:19]
  wire  m_914_io_s; // @[MUL.scala 102:19]
  wire  m_914_io_cout; // @[MUL.scala 102:19]
  wire  m_915_io_x1; // @[MUL.scala 102:19]
  wire  m_915_io_x2; // @[MUL.scala 102:19]
  wire  m_915_io_x3; // @[MUL.scala 102:19]
  wire  m_915_io_s; // @[MUL.scala 102:19]
  wire  m_915_io_cout; // @[MUL.scala 102:19]
  wire  m_916_io_x1; // @[MUL.scala 102:19]
  wire  m_916_io_x2; // @[MUL.scala 102:19]
  wire  m_916_io_x3; // @[MUL.scala 102:19]
  wire  m_916_io_s; // @[MUL.scala 102:19]
  wire  m_916_io_cout; // @[MUL.scala 102:19]
  wire  m_917_io_x1; // @[MUL.scala 102:19]
  wire  m_917_io_x2; // @[MUL.scala 102:19]
  wire  m_917_io_x3; // @[MUL.scala 102:19]
  wire  m_917_io_s; // @[MUL.scala 102:19]
  wire  m_917_io_cout; // @[MUL.scala 102:19]
  wire  m_918_io_x1; // @[MUL.scala 102:19]
  wire  m_918_io_x2; // @[MUL.scala 102:19]
  wire  m_918_io_x3; // @[MUL.scala 102:19]
  wire  m_918_io_s; // @[MUL.scala 102:19]
  wire  m_918_io_cout; // @[MUL.scala 102:19]
  wire  m_919_io_x1; // @[MUL.scala 102:19]
  wire  m_919_io_x2; // @[MUL.scala 102:19]
  wire  m_919_io_x3; // @[MUL.scala 102:19]
  wire  m_919_io_s; // @[MUL.scala 102:19]
  wire  m_919_io_cout; // @[MUL.scala 102:19]
  wire  m_920_io_x1; // @[MUL.scala 102:19]
  wire  m_920_io_x2; // @[MUL.scala 102:19]
  wire  m_920_io_x3; // @[MUL.scala 102:19]
  wire  m_920_io_s; // @[MUL.scala 102:19]
  wire  m_920_io_cout; // @[MUL.scala 102:19]
  wire  m_921_io_x1; // @[MUL.scala 102:19]
  wire  m_921_io_x2; // @[MUL.scala 102:19]
  wire  m_921_io_x3; // @[MUL.scala 102:19]
  wire  m_921_io_s; // @[MUL.scala 102:19]
  wire  m_921_io_cout; // @[MUL.scala 102:19]
  wire  m_922_io_x1; // @[MUL.scala 102:19]
  wire  m_922_io_x2; // @[MUL.scala 102:19]
  wire  m_922_io_x3; // @[MUL.scala 102:19]
  wire  m_922_io_s; // @[MUL.scala 102:19]
  wire  m_922_io_cout; // @[MUL.scala 102:19]
  wire  m_923_io_x1; // @[MUL.scala 102:19]
  wire  m_923_io_x2; // @[MUL.scala 102:19]
  wire  m_923_io_x3; // @[MUL.scala 102:19]
  wire  m_923_io_s; // @[MUL.scala 102:19]
  wire  m_923_io_cout; // @[MUL.scala 102:19]
  wire  m_924_io_x1; // @[MUL.scala 102:19]
  wire  m_924_io_x2; // @[MUL.scala 102:19]
  wire  m_924_io_x3; // @[MUL.scala 102:19]
  wire  m_924_io_s; // @[MUL.scala 102:19]
  wire  m_924_io_cout; // @[MUL.scala 102:19]
  wire  m_925_io_x1; // @[MUL.scala 102:19]
  wire  m_925_io_x2; // @[MUL.scala 102:19]
  wire  m_925_io_x3; // @[MUL.scala 102:19]
  wire  m_925_io_s; // @[MUL.scala 102:19]
  wire  m_925_io_cout; // @[MUL.scala 102:19]
  wire  m_926_io_x1; // @[MUL.scala 102:19]
  wire  m_926_io_x2; // @[MUL.scala 102:19]
  wire  m_926_io_x3; // @[MUL.scala 102:19]
  wire  m_926_io_s; // @[MUL.scala 102:19]
  wire  m_926_io_cout; // @[MUL.scala 102:19]
  wire  m_927_io_x1; // @[MUL.scala 102:19]
  wire  m_927_io_x2; // @[MUL.scala 102:19]
  wire  m_927_io_x3; // @[MUL.scala 102:19]
  wire  m_927_io_s; // @[MUL.scala 102:19]
  wire  m_927_io_cout; // @[MUL.scala 102:19]
  wire  m_928_io_x1; // @[MUL.scala 102:19]
  wire  m_928_io_x2; // @[MUL.scala 102:19]
  wire  m_928_io_x3; // @[MUL.scala 102:19]
  wire  m_928_io_s; // @[MUL.scala 102:19]
  wire  m_928_io_cout; // @[MUL.scala 102:19]
  wire  m_929_io_x1; // @[MUL.scala 102:19]
  wire  m_929_io_x2; // @[MUL.scala 102:19]
  wire  m_929_io_x3; // @[MUL.scala 102:19]
  wire  m_929_io_s; // @[MUL.scala 102:19]
  wire  m_929_io_cout; // @[MUL.scala 102:19]
  wire  m_930_io_x1; // @[MUL.scala 102:19]
  wire  m_930_io_x2; // @[MUL.scala 102:19]
  wire  m_930_io_x3; // @[MUL.scala 102:19]
  wire  m_930_io_s; // @[MUL.scala 102:19]
  wire  m_930_io_cout; // @[MUL.scala 102:19]
  wire  m_931_io_x1; // @[MUL.scala 102:19]
  wire  m_931_io_x2; // @[MUL.scala 102:19]
  wire  m_931_io_x3; // @[MUL.scala 102:19]
  wire  m_931_io_s; // @[MUL.scala 102:19]
  wire  m_931_io_cout; // @[MUL.scala 102:19]
  wire  m_932_io_x1; // @[MUL.scala 102:19]
  wire  m_932_io_x2; // @[MUL.scala 102:19]
  wire  m_932_io_x3; // @[MUL.scala 102:19]
  wire  m_932_io_s; // @[MUL.scala 102:19]
  wire  m_932_io_cout; // @[MUL.scala 102:19]
  wire  m_933_io_x1; // @[MUL.scala 102:19]
  wire  m_933_io_x2; // @[MUL.scala 102:19]
  wire  m_933_io_x3; // @[MUL.scala 102:19]
  wire  m_933_io_s; // @[MUL.scala 102:19]
  wire  m_933_io_cout; // @[MUL.scala 102:19]
  wire  m_934_io_x1; // @[MUL.scala 102:19]
  wire  m_934_io_x2; // @[MUL.scala 102:19]
  wire  m_934_io_x3; // @[MUL.scala 102:19]
  wire  m_934_io_s; // @[MUL.scala 102:19]
  wire  m_934_io_cout; // @[MUL.scala 102:19]
  wire  m_935_io_x1; // @[MUL.scala 102:19]
  wire  m_935_io_x2; // @[MUL.scala 102:19]
  wire  m_935_io_x3; // @[MUL.scala 102:19]
  wire  m_935_io_s; // @[MUL.scala 102:19]
  wire  m_935_io_cout; // @[MUL.scala 102:19]
  wire  m_936_io_x1; // @[MUL.scala 102:19]
  wire  m_936_io_x2; // @[MUL.scala 102:19]
  wire  m_936_io_x3; // @[MUL.scala 102:19]
  wire  m_936_io_s; // @[MUL.scala 102:19]
  wire  m_936_io_cout; // @[MUL.scala 102:19]
  wire  m_937_io_x1; // @[MUL.scala 102:19]
  wire  m_937_io_x2; // @[MUL.scala 102:19]
  wire  m_937_io_x3; // @[MUL.scala 102:19]
  wire  m_937_io_s; // @[MUL.scala 102:19]
  wire  m_937_io_cout; // @[MUL.scala 102:19]
  wire  m_938_io_x1; // @[MUL.scala 102:19]
  wire  m_938_io_x2; // @[MUL.scala 102:19]
  wire  m_938_io_x3; // @[MUL.scala 102:19]
  wire  m_938_io_s; // @[MUL.scala 102:19]
  wire  m_938_io_cout; // @[MUL.scala 102:19]
  wire  m_939_io_x1; // @[MUL.scala 102:19]
  wire  m_939_io_x2; // @[MUL.scala 102:19]
  wire  m_939_io_x3; // @[MUL.scala 102:19]
  wire  m_939_io_s; // @[MUL.scala 102:19]
  wire  m_939_io_cout; // @[MUL.scala 102:19]
  wire  m_940_io_x1; // @[MUL.scala 102:19]
  wire  m_940_io_x2; // @[MUL.scala 102:19]
  wire  m_940_io_x3; // @[MUL.scala 102:19]
  wire  m_940_io_s; // @[MUL.scala 102:19]
  wire  m_940_io_cout; // @[MUL.scala 102:19]
  wire  m_941_io_x1; // @[MUL.scala 102:19]
  wire  m_941_io_x2; // @[MUL.scala 102:19]
  wire  m_941_io_x3; // @[MUL.scala 102:19]
  wire  m_941_io_s; // @[MUL.scala 102:19]
  wire  m_941_io_cout; // @[MUL.scala 102:19]
  wire  m_942_io_x1; // @[MUL.scala 102:19]
  wire  m_942_io_x2; // @[MUL.scala 102:19]
  wire  m_942_io_x3; // @[MUL.scala 102:19]
  wire  m_942_io_s; // @[MUL.scala 102:19]
  wire  m_942_io_cout; // @[MUL.scala 102:19]
  wire  m_943_io_in_0; // @[MUL.scala 124:19]
  wire  m_943_io_in_1; // @[MUL.scala 124:19]
  wire  m_943_io_out_0; // @[MUL.scala 124:19]
  wire  m_943_io_out_1; // @[MUL.scala 124:19]
  wire  m_944_io_x1; // @[MUL.scala 102:19]
  wire  m_944_io_x2; // @[MUL.scala 102:19]
  wire  m_944_io_x3; // @[MUL.scala 102:19]
  wire  m_944_io_s; // @[MUL.scala 102:19]
  wire  m_944_io_cout; // @[MUL.scala 102:19]
  wire  m_945_io_x1; // @[MUL.scala 102:19]
  wire  m_945_io_x2; // @[MUL.scala 102:19]
  wire  m_945_io_x3; // @[MUL.scala 102:19]
  wire  m_945_io_s; // @[MUL.scala 102:19]
  wire  m_945_io_cout; // @[MUL.scala 102:19]
  wire  m_946_io_x1; // @[MUL.scala 102:19]
  wire  m_946_io_x2; // @[MUL.scala 102:19]
  wire  m_946_io_x3; // @[MUL.scala 102:19]
  wire  m_946_io_s; // @[MUL.scala 102:19]
  wire  m_946_io_cout; // @[MUL.scala 102:19]
  wire  m_947_io_x1; // @[MUL.scala 102:19]
  wire  m_947_io_x2; // @[MUL.scala 102:19]
  wire  m_947_io_x3; // @[MUL.scala 102:19]
  wire  m_947_io_s; // @[MUL.scala 102:19]
  wire  m_947_io_cout; // @[MUL.scala 102:19]
  wire  m_948_io_x1; // @[MUL.scala 102:19]
  wire  m_948_io_x2; // @[MUL.scala 102:19]
  wire  m_948_io_x3; // @[MUL.scala 102:19]
  wire  m_948_io_s; // @[MUL.scala 102:19]
  wire  m_948_io_cout; // @[MUL.scala 102:19]
  wire  m_949_io_in_0; // @[MUL.scala 124:19]
  wire  m_949_io_in_1; // @[MUL.scala 124:19]
  wire  m_949_io_out_0; // @[MUL.scala 124:19]
  wire  m_949_io_out_1; // @[MUL.scala 124:19]
  wire  m_950_io_x1; // @[MUL.scala 102:19]
  wire  m_950_io_x2; // @[MUL.scala 102:19]
  wire  m_950_io_x3; // @[MUL.scala 102:19]
  wire  m_950_io_s; // @[MUL.scala 102:19]
  wire  m_950_io_cout; // @[MUL.scala 102:19]
  wire  m_951_io_x1; // @[MUL.scala 102:19]
  wire  m_951_io_x2; // @[MUL.scala 102:19]
  wire  m_951_io_x3; // @[MUL.scala 102:19]
  wire  m_951_io_s; // @[MUL.scala 102:19]
  wire  m_951_io_cout; // @[MUL.scala 102:19]
  wire  m_952_io_x1; // @[MUL.scala 102:19]
  wire  m_952_io_x2; // @[MUL.scala 102:19]
  wire  m_952_io_x3; // @[MUL.scala 102:19]
  wire  m_952_io_s; // @[MUL.scala 102:19]
  wire  m_952_io_cout; // @[MUL.scala 102:19]
  wire  m_953_io_x1; // @[MUL.scala 102:19]
  wire  m_953_io_x2; // @[MUL.scala 102:19]
  wire  m_953_io_x3; // @[MUL.scala 102:19]
  wire  m_953_io_s; // @[MUL.scala 102:19]
  wire  m_953_io_cout; // @[MUL.scala 102:19]
  wire  m_954_io_x1; // @[MUL.scala 102:19]
  wire  m_954_io_x2; // @[MUL.scala 102:19]
  wire  m_954_io_x3; // @[MUL.scala 102:19]
  wire  m_954_io_s; // @[MUL.scala 102:19]
  wire  m_954_io_cout; // @[MUL.scala 102:19]
  wire  m_955_io_in_0; // @[MUL.scala 124:19]
  wire  m_955_io_in_1; // @[MUL.scala 124:19]
  wire  m_955_io_out_0; // @[MUL.scala 124:19]
  wire  m_955_io_out_1; // @[MUL.scala 124:19]
  wire  m_956_io_x1; // @[MUL.scala 102:19]
  wire  m_956_io_x2; // @[MUL.scala 102:19]
  wire  m_956_io_x3; // @[MUL.scala 102:19]
  wire  m_956_io_s; // @[MUL.scala 102:19]
  wire  m_956_io_cout; // @[MUL.scala 102:19]
  wire  m_957_io_x1; // @[MUL.scala 102:19]
  wire  m_957_io_x2; // @[MUL.scala 102:19]
  wire  m_957_io_x3; // @[MUL.scala 102:19]
  wire  m_957_io_s; // @[MUL.scala 102:19]
  wire  m_957_io_cout; // @[MUL.scala 102:19]
  wire  m_958_io_x1; // @[MUL.scala 102:19]
  wire  m_958_io_x2; // @[MUL.scala 102:19]
  wire  m_958_io_x3; // @[MUL.scala 102:19]
  wire  m_958_io_s; // @[MUL.scala 102:19]
  wire  m_958_io_cout; // @[MUL.scala 102:19]
  wire  m_959_io_x1; // @[MUL.scala 102:19]
  wire  m_959_io_x2; // @[MUL.scala 102:19]
  wire  m_959_io_x3; // @[MUL.scala 102:19]
  wire  m_959_io_s; // @[MUL.scala 102:19]
  wire  m_959_io_cout; // @[MUL.scala 102:19]
  wire  m_960_io_x1; // @[MUL.scala 102:19]
  wire  m_960_io_x2; // @[MUL.scala 102:19]
  wire  m_960_io_x3; // @[MUL.scala 102:19]
  wire  m_960_io_s; // @[MUL.scala 102:19]
  wire  m_960_io_cout; // @[MUL.scala 102:19]
  wire  m_961_io_x1; // @[MUL.scala 102:19]
  wire  m_961_io_x2; // @[MUL.scala 102:19]
  wire  m_961_io_x3; // @[MUL.scala 102:19]
  wire  m_961_io_s; // @[MUL.scala 102:19]
  wire  m_961_io_cout; // @[MUL.scala 102:19]
  wire  m_962_io_x1; // @[MUL.scala 102:19]
  wire  m_962_io_x2; // @[MUL.scala 102:19]
  wire  m_962_io_x3; // @[MUL.scala 102:19]
  wire  m_962_io_s; // @[MUL.scala 102:19]
  wire  m_962_io_cout; // @[MUL.scala 102:19]
  wire  m_963_io_x1; // @[MUL.scala 102:19]
  wire  m_963_io_x2; // @[MUL.scala 102:19]
  wire  m_963_io_x3; // @[MUL.scala 102:19]
  wire  m_963_io_s; // @[MUL.scala 102:19]
  wire  m_963_io_cout; // @[MUL.scala 102:19]
  wire  m_964_io_x1; // @[MUL.scala 102:19]
  wire  m_964_io_x2; // @[MUL.scala 102:19]
  wire  m_964_io_x3; // @[MUL.scala 102:19]
  wire  m_964_io_s; // @[MUL.scala 102:19]
  wire  m_964_io_cout; // @[MUL.scala 102:19]
  wire  m_965_io_x1; // @[MUL.scala 102:19]
  wire  m_965_io_x2; // @[MUL.scala 102:19]
  wire  m_965_io_x3; // @[MUL.scala 102:19]
  wire  m_965_io_s; // @[MUL.scala 102:19]
  wire  m_965_io_cout; // @[MUL.scala 102:19]
  wire  m_966_io_x1; // @[MUL.scala 102:19]
  wire  m_966_io_x2; // @[MUL.scala 102:19]
  wire  m_966_io_x3; // @[MUL.scala 102:19]
  wire  m_966_io_s; // @[MUL.scala 102:19]
  wire  m_966_io_cout; // @[MUL.scala 102:19]
  wire  m_967_io_x1; // @[MUL.scala 102:19]
  wire  m_967_io_x2; // @[MUL.scala 102:19]
  wire  m_967_io_x3; // @[MUL.scala 102:19]
  wire  m_967_io_s; // @[MUL.scala 102:19]
  wire  m_967_io_cout; // @[MUL.scala 102:19]
  wire  m_968_io_x1; // @[MUL.scala 102:19]
  wire  m_968_io_x2; // @[MUL.scala 102:19]
  wire  m_968_io_x3; // @[MUL.scala 102:19]
  wire  m_968_io_s; // @[MUL.scala 102:19]
  wire  m_968_io_cout; // @[MUL.scala 102:19]
  wire  m_969_io_x1; // @[MUL.scala 102:19]
  wire  m_969_io_x2; // @[MUL.scala 102:19]
  wire  m_969_io_x3; // @[MUL.scala 102:19]
  wire  m_969_io_s; // @[MUL.scala 102:19]
  wire  m_969_io_cout; // @[MUL.scala 102:19]
  wire  m_970_io_x1; // @[MUL.scala 102:19]
  wire  m_970_io_x2; // @[MUL.scala 102:19]
  wire  m_970_io_x3; // @[MUL.scala 102:19]
  wire  m_970_io_s; // @[MUL.scala 102:19]
  wire  m_970_io_cout; // @[MUL.scala 102:19]
  wire  m_971_io_x1; // @[MUL.scala 102:19]
  wire  m_971_io_x2; // @[MUL.scala 102:19]
  wire  m_971_io_x3; // @[MUL.scala 102:19]
  wire  m_971_io_s; // @[MUL.scala 102:19]
  wire  m_971_io_cout; // @[MUL.scala 102:19]
  wire  m_972_io_x1; // @[MUL.scala 102:19]
  wire  m_972_io_x2; // @[MUL.scala 102:19]
  wire  m_972_io_x3; // @[MUL.scala 102:19]
  wire  m_972_io_s; // @[MUL.scala 102:19]
  wire  m_972_io_cout; // @[MUL.scala 102:19]
  wire  m_973_io_x1; // @[MUL.scala 102:19]
  wire  m_973_io_x2; // @[MUL.scala 102:19]
  wire  m_973_io_x3; // @[MUL.scala 102:19]
  wire  m_973_io_s; // @[MUL.scala 102:19]
  wire  m_973_io_cout; // @[MUL.scala 102:19]
  wire  m_974_io_x1; // @[MUL.scala 102:19]
  wire  m_974_io_x2; // @[MUL.scala 102:19]
  wire  m_974_io_x3; // @[MUL.scala 102:19]
  wire  m_974_io_s; // @[MUL.scala 102:19]
  wire  m_974_io_cout; // @[MUL.scala 102:19]
  wire  m_975_io_x1; // @[MUL.scala 102:19]
  wire  m_975_io_x2; // @[MUL.scala 102:19]
  wire  m_975_io_x3; // @[MUL.scala 102:19]
  wire  m_975_io_s; // @[MUL.scala 102:19]
  wire  m_975_io_cout; // @[MUL.scala 102:19]
  wire  m_976_io_x1; // @[MUL.scala 102:19]
  wire  m_976_io_x2; // @[MUL.scala 102:19]
  wire  m_976_io_x3; // @[MUL.scala 102:19]
  wire  m_976_io_s; // @[MUL.scala 102:19]
  wire  m_976_io_cout; // @[MUL.scala 102:19]
  wire  m_977_io_x1; // @[MUL.scala 102:19]
  wire  m_977_io_x2; // @[MUL.scala 102:19]
  wire  m_977_io_x3; // @[MUL.scala 102:19]
  wire  m_977_io_s; // @[MUL.scala 102:19]
  wire  m_977_io_cout; // @[MUL.scala 102:19]
  wire  m_978_io_x1; // @[MUL.scala 102:19]
  wire  m_978_io_x2; // @[MUL.scala 102:19]
  wire  m_978_io_x3; // @[MUL.scala 102:19]
  wire  m_978_io_s; // @[MUL.scala 102:19]
  wire  m_978_io_cout; // @[MUL.scala 102:19]
  wire  m_979_io_x1; // @[MUL.scala 102:19]
  wire  m_979_io_x2; // @[MUL.scala 102:19]
  wire  m_979_io_x3; // @[MUL.scala 102:19]
  wire  m_979_io_s; // @[MUL.scala 102:19]
  wire  m_979_io_cout; // @[MUL.scala 102:19]
  wire  m_980_io_x1; // @[MUL.scala 102:19]
  wire  m_980_io_x2; // @[MUL.scala 102:19]
  wire  m_980_io_x3; // @[MUL.scala 102:19]
  wire  m_980_io_s; // @[MUL.scala 102:19]
  wire  m_980_io_cout; // @[MUL.scala 102:19]
  wire  m_981_io_x1; // @[MUL.scala 102:19]
  wire  m_981_io_x2; // @[MUL.scala 102:19]
  wire  m_981_io_x3; // @[MUL.scala 102:19]
  wire  m_981_io_s; // @[MUL.scala 102:19]
  wire  m_981_io_cout; // @[MUL.scala 102:19]
  wire  m_982_io_x1; // @[MUL.scala 102:19]
  wire  m_982_io_x2; // @[MUL.scala 102:19]
  wire  m_982_io_x3; // @[MUL.scala 102:19]
  wire  m_982_io_s; // @[MUL.scala 102:19]
  wire  m_982_io_cout; // @[MUL.scala 102:19]
  wire  m_983_io_x1; // @[MUL.scala 102:19]
  wire  m_983_io_x2; // @[MUL.scala 102:19]
  wire  m_983_io_x3; // @[MUL.scala 102:19]
  wire  m_983_io_s; // @[MUL.scala 102:19]
  wire  m_983_io_cout; // @[MUL.scala 102:19]
  wire  m_984_io_x1; // @[MUL.scala 102:19]
  wire  m_984_io_x2; // @[MUL.scala 102:19]
  wire  m_984_io_x3; // @[MUL.scala 102:19]
  wire  m_984_io_s; // @[MUL.scala 102:19]
  wire  m_984_io_cout; // @[MUL.scala 102:19]
  wire  m_985_io_x1; // @[MUL.scala 102:19]
  wire  m_985_io_x2; // @[MUL.scala 102:19]
  wire  m_985_io_x3; // @[MUL.scala 102:19]
  wire  m_985_io_s; // @[MUL.scala 102:19]
  wire  m_985_io_cout; // @[MUL.scala 102:19]
  wire  m_986_io_x1; // @[MUL.scala 102:19]
  wire  m_986_io_x2; // @[MUL.scala 102:19]
  wire  m_986_io_x3; // @[MUL.scala 102:19]
  wire  m_986_io_s; // @[MUL.scala 102:19]
  wire  m_986_io_cout; // @[MUL.scala 102:19]
  wire  m_987_io_x1; // @[MUL.scala 102:19]
  wire  m_987_io_x2; // @[MUL.scala 102:19]
  wire  m_987_io_x3; // @[MUL.scala 102:19]
  wire  m_987_io_s; // @[MUL.scala 102:19]
  wire  m_987_io_cout; // @[MUL.scala 102:19]
  wire  m_988_io_x1; // @[MUL.scala 102:19]
  wire  m_988_io_x2; // @[MUL.scala 102:19]
  wire  m_988_io_x3; // @[MUL.scala 102:19]
  wire  m_988_io_s; // @[MUL.scala 102:19]
  wire  m_988_io_cout; // @[MUL.scala 102:19]
  wire  m_989_io_x1; // @[MUL.scala 102:19]
  wire  m_989_io_x2; // @[MUL.scala 102:19]
  wire  m_989_io_x3; // @[MUL.scala 102:19]
  wire  m_989_io_s; // @[MUL.scala 102:19]
  wire  m_989_io_cout; // @[MUL.scala 102:19]
  wire  m_990_io_x1; // @[MUL.scala 102:19]
  wire  m_990_io_x2; // @[MUL.scala 102:19]
  wire  m_990_io_x3; // @[MUL.scala 102:19]
  wire  m_990_io_s; // @[MUL.scala 102:19]
  wire  m_990_io_cout; // @[MUL.scala 102:19]
  wire  m_991_io_x1; // @[MUL.scala 102:19]
  wire  m_991_io_x2; // @[MUL.scala 102:19]
  wire  m_991_io_x3; // @[MUL.scala 102:19]
  wire  m_991_io_s; // @[MUL.scala 102:19]
  wire  m_991_io_cout; // @[MUL.scala 102:19]
  wire  m_992_io_x1; // @[MUL.scala 102:19]
  wire  m_992_io_x2; // @[MUL.scala 102:19]
  wire  m_992_io_x3; // @[MUL.scala 102:19]
  wire  m_992_io_s; // @[MUL.scala 102:19]
  wire  m_992_io_cout; // @[MUL.scala 102:19]
  wire  m_993_io_x1; // @[MUL.scala 102:19]
  wire  m_993_io_x2; // @[MUL.scala 102:19]
  wire  m_993_io_x3; // @[MUL.scala 102:19]
  wire  m_993_io_s; // @[MUL.scala 102:19]
  wire  m_993_io_cout; // @[MUL.scala 102:19]
  wire  m_994_io_x1; // @[MUL.scala 102:19]
  wire  m_994_io_x2; // @[MUL.scala 102:19]
  wire  m_994_io_x3; // @[MUL.scala 102:19]
  wire  m_994_io_s; // @[MUL.scala 102:19]
  wire  m_994_io_cout; // @[MUL.scala 102:19]
  wire  m_995_io_x1; // @[MUL.scala 102:19]
  wire  m_995_io_x2; // @[MUL.scala 102:19]
  wire  m_995_io_x3; // @[MUL.scala 102:19]
  wire  m_995_io_s; // @[MUL.scala 102:19]
  wire  m_995_io_cout; // @[MUL.scala 102:19]
  wire  m_996_io_x1; // @[MUL.scala 102:19]
  wire  m_996_io_x2; // @[MUL.scala 102:19]
  wire  m_996_io_x3; // @[MUL.scala 102:19]
  wire  m_996_io_s; // @[MUL.scala 102:19]
  wire  m_996_io_cout; // @[MUL.scala 102:19]
  wire  m_997_io_x1; // @[MUL.scala 102:19]
  wire  m_997_io_x2; // @[MUL.scala 102:19]
  wire  m_997_io_x3; // @[MUL.scala 102:19]
  wire  m_997_io_s; // @[MUL.scala 102:19]
  wire  m_997_io_cout; // @[MUL.scala 102:19]
  wire  m_998_io_in_0; // @[MUL.scala 124:19]
  wire  m_998_io_in_1; // @[MUL.scala 124:19]
  wire  m_998_io_out_0; // @[MUL.scala 124:19]
  wire  m_998_io_out_1; // @[MUL.scala 124:19]
  wire  m_999_io_x1; // @[MUL.scala 102:19]
  wire  m_999_io_x2; // @[MUL.scala 102:19]
  wire  m_999_io_x3; // @[MUL.scala 102:19]
  wire  m_999_io_s; // @[MUL.scala 102:19]
  wire  m_999_io_cout; // @[MUL.scala 102:19]
  wire  m_1000_io_x1; // @[MUL.scala 102:19]
  wire  m_1000_io_x2; // @[MUL.scala 102:19]
  wire  m_1000_io_x3; // @[MUL.scala 102:19]
  wire  m_1000_io_s; // @[MUL.scala 102:19]
  wire  m_1000_io_cout; // @[MUL.scala 102:19]
  wire  m_1001_io_x1; // @[MUL.scala 102:19]
  wire  m_1001_io_x2; // @[MUL.scala 102:19]
  wire  m_1001_io_x3; // @[MUL.scala 102:19]
  wire  m_1001_io_s; // @[MUL.scala 102:19]
  wire  m_1001_io_cout; // @[MUL.scala 102:19]
  wire  m_1002_io_x1; // @[MUL.scala 102:19]
  wire  m_1002_io_x2; // @[MUL.scala 102:19]
  wire  m_1002_io_x3; // @[MUL.scala 102:19]
  wire  m_1002_io_s; // @[MUL.scala 102:19]
  wire  m_1002_io_cout; // @[MUL.scala 102:19]
  wire  m_1003_io_x1; // @[MUL.scala 102:19]
  wire  m_1003_io_x2; // @[MUL.scala 102:19]
  wire  m_1003_io_x3; // @[MUL.scala 102:19]
  wire  m_1003_io_s; // @[MUL.scala 102:19]
  wire  m_1003_io_cout; // @[MUL.scala 102:19]
  wire  m_1004_io_x1; // @[MUL.scala 102:19]
  wire  m_1004_io_x2; // @[MUL.scala 102:19]
  wire  m_1004_io_x3; // @[MUL.scala 102:19]
  wire  m_1004_io_s; // @[MUL.scala 102:19]
  wire  m_1004_io_cout; // @[MUL.scala 102:19]
  wire  m_1005_io_in_0; // @[MUL.scala 124:19]
  wire  m_1005_io_in_1; // @[MUL.scala 124:19]
  wire  m_1005_io_out_0; // @[MUL.scala 124:19]
  wire  m_1005_io_out_1; // @[MUL.scala 124:19]
  wire  m_1006_io_x1; // @[MUL.scala 102:19]
  wire  m_1006_io_x2; // @[MUL.scala 102:19]
  wire  m_1006_io_x3; // @[MUL.scala 102:19]
  wire  m_1006_io_s; // @[MUL.scala 102:19]
  wire  m_1006_io_cout; // @[MUL.scala 102:19]
  wire  m_1007_io_x1; // @[MUL.scala 102:19]
  wire  m_1007_io_x2; // @[MUL.scala 102:19]
  wire  m_1007_io_x3; // @[MUL.scala 102:19]
  wire  m_1007_io_s; // @[MUL.scala 102:19]
  wire  m_1007_io_cout; // @[MUL.scala 102:19]
  wire  m_1008_io_x1; // @[MUL.scala 102:19]
  wire  m_1008_io_x2; // @[MUL.scala 102:19]
  wire  m_1008_io_x3; // @[MUL.scala 102:19]
  wire  m_1008_io_s; // @[MUL.scala 102:19]
  wire  m_1008_io_cout; // @[MUL.scala 102:19]
  wire  m_1009_io_x1; // @[MUL.scala 102:19]
  wire  m_1009_io_x2; // @[MUL.scala 102:19]
  wire  m_1009_io_x3; // @[MUL.scala 102:19]
  wire  m_1009_io_s; // @[MUL.scala 102:19]
  wire  m_1009_io_cout; // @[MUL.scala 102:19]
  wire  m_1010_io_x1; // @[MUL.scala 102:19]
  wire  m_1010_io_x2; // @[MUL.scala 102:19]
  wire  m_1010_io_x3; // @[MUL.scala 102:19]
  wire  m_1010_io_s; // @[MUL.scala 102:19]
  wire  m_1010_io_cout; // @[MUL.scala 102:19]
  wire  m_1011_io_x1; // @[MUL.scala 102:19]
  wire  m_1011_io_x2; // @[MUL.scala 102:19]
  wire  m_1011_io_x3; // @[MUL.scala 102:19]
  wire  m_1011_io_s; // @[MUL.scala 102:19]
  wire  m_1011_io_cout; // @[MUL.scala 102:19]
  wire  m_1012_io_in_0; // @[MUL.scala 124:19]
  wire  m_1012_io_in_1; // @[MUL.scala 124:19]
  wire  m_1012_io_out_0; // @[MUL.scala 124:19]
  wire  m_1012_io_out_1; // @[MUL.scala 124:19]
  wire  m_1013_io_x1; // @[MUL.scala 102:19]
  wire  m_1013_io_x2; // @[MUL.scala 102:19]
  wire  m_1013_io_x3; // @[MUL.scala 102:19]
  wire  m_1013_io_s; // @[MUL.scala 102:19]
  wire  m_1013_io_cout; // @[MUL.scala 102:19]
  wire  m_1014_io_x1; // @[MUL.scala 102:19]
  wire  m_1014_io_x2; // @[MUL.scala 102:19]
  wire  m_1014_io_x3; // @[MUL.scala 102:19]
  wire  m_1014_io_s; // @[MUL.scala 102:19]
  wire  m_1014_io_cout; // @[MUL.scala 102:19]
  wire  m_1015_io_x1; // @[MUL.scala 102:19]
  wire  m_1015_io_x2; // @[MUL.scala 102:19]
  wire  m_1015_io_x3; // @[MUL.scala 102:19]
  wire  m_1015_io_s; // @[MUL.scala 102:19]
  wire  m_1015_io_cout; // @[MUL.scala 102:19]
  wire  m_1016_io_x1; // @[MUL.scala 102:19]
  wire  m_1016_io_x2; // @[MUL.scala 102:19]
  wire  m_1016_io_x3; // @[MUL.scala 102:19]
  wire  m_1016_io_s; // @[MUL.scala 102:19]
  wire  m_1016_io_cout; // @[MUL.scala 102:19]
  wire  m_1017_io_x1; // @[MUL.scala 102:19]
  wire  m_1017_io_x2; // @[MUL.scala 102:19]
  wire  m_1017_io_x3; // @[MUL.scala 102:19]
  wire  m_1017_io_s; // @[MUL.scala 102:19]
  wire  m_1017_io_cout; // @[MUL.scala 102:19]
  wire  m_1018_io_x1; // @[MUL.scala 102:19]
  wire  m_1018_io_x2; // @[MUL.scala 102:19]
  wire  m_1018_io_x3; // @[MUL.scala 102:19]
  wire  m_1018_io_s; // @[MUL.scala 102:19]
  wire  m_1018_io_cout; // @[MUL.scala 102:19]
  wire  m_1019_io_x1; // @[MUL.scala 102:19]
  wire  m_1019_io_x2; // @[MUL.scala 102:19]
  wire  m_1019_io_x3; // @[MUL.scala 102:19]
  wire  m_1019_io_s; // @[MUL.scala 102:19]
  wire  m_1019_io_cout; // @[MUL.scala 102:19]
  wire  m_1020_io_x1; // @[MUL.scala 102:19]
  wire  m_1020_io_x2; // @[MUL.scala 102:19]
  wire  m_1020_io_x3; // @[MUL.scala 102:19]
  wire  m_1020_io_s; // @[MUL.scala 102:19]
  wire  m_1020_io_cout; // @[MUL.scala 102:19]
  wire  m_1021_io_x1; // @[MUL.scala 102:19]
  wire  m_1021_io_x2; // @[MUL.scala 102:19]
  wire  m_1021_io_x3; // @[MUL.scala 102:19]
  wire  m_1021_io_s; // @[MUL.scala 102:19]
  wire  m_1021_io_cout; // @[MUL.scala 102:19]
  wire  m_1022_io_x1; // @[MUL.scala 102:19]
  wire  m_1022_io_x2; // @[MUL.scala 102:19]
  wire  m_1022_io_x3; // @[MUL.scala 102:19]
  wire  m_1022_io_s; // @[MUL.scala 102:19]
  wire  m_1022_io_cout; // @[MUL.scala 102:19]
  wire  m_1023_io_x1; // @[MUL.scala 102:19]
  wire  m_1023_io_x2; // @[MUL.scala 102:19]
  wire  m_1023_io_x3; // @[MUL.scala 102:19]
  wire  m_1023_io_s; // @[MUL.scala 102:19]
  wire  m_1023_io_cout; // @[MUL.scala 102:19]
  wire  m_1024_io_x1; // @[MUL.scala 102:19]
  wire  m_1024_io_x2; // @[MUL.scala 102:19]
  wire  m_1024_io_x3; // @[MUL.scala 102:19]
  wire  m_1024_io_s; // @[MUL.scala 102:19]
  wire  m_1024_io_cout; // @[MUL.scala 102:19]
  wire  m_1025_io_x1; // @[MUL.scala 102:19]
  wire  m_1025_io_x2; // @[MUL.scala 102:19]
  wire  m_1025_io_x3; // @[MUL.scala 102:19]
  wire  m_1025_io_s; // @[MUL.scala 102:19]
  wire  m_1025_io_cout; // @[MUL.scala 102:19]
  wire  m_1026_io_x1; // @[MUL.scala 102:19]
  wire  m_1026_io_x2; // @[MUL.scala 102:19]
  wire  m_1026_io_x3; // @[MUL.scala 102:19]
  wire  m_1026_io_s; // @[MUL.scala 102:19]
  wire  m_1026_io_cout; // @[MUL.scala 102:19]
  wire  m_1027_io_x1; // @[MUL.scala 102:19]
  wire  m_1027_io_x2; // @[MUL.scala 102:19]
  wire  m_1027_io_x3; // @[MUL.scala 102:19]
  wire  m_1027_io_s; // @[MUL.scala 102:19]
  wire  m_1027_io_cout; // @[MUL.scala 102:19]
  wire  m_1028_io_x1; // @[MUL.scala 102:19]
  wire  m_1028_io_x2; // @[MUL.scala 102:19]
  wire  m_1028_io_x3; // @[MUL.scala 102:19]
  wire  m_1028_io_s; // @[MUL.scala 102:19]
  wire  m_1028_io_cout; // @[MUL.scala 102:19]
  wire  m_1029_io_x1; // @[MUL.scala 102:19]
  wire  m_1029_io_x2; // @[MUL.scala 102:19]
  wire  m_1029_io_x3; // @[MUL.scala 102:19]
  wire  m_1029_io_s; // @[MUL.scala 102:19]
  wire  m_1029_io_cout; // @[MUL.scala 102:19]
  wire  m_1030_io_x1; // @[MUL.scala 102:19]
  wire  m_1030_io_x2; // @[MUL.scala 102:19]
  wire  m_1030_io_x3; // @[MUL.scala 102:19]
  wire  m_1030_io_s; // @[MUL.scala 102:19]
  wire  m_1030_io_cout; // @[MUL.scala 102:19]
  wire  m_1031_io_x1; // @[MUL.scala 102:19]
  wire  m_1031_io_x2; // @[MUL.scala 102:19]
  wire  m_1031_io_x3; // @[MUL.scala 102:19]
  wire  m_1031_io_s; // @[MUL.scala 102:19]
  wire  m_1031_io_cout; // @[MUL.scala 102:19]
  wire  m_1032_io_x1; // @[MUL.scala 102:19]
  wire  m_1032_io_x2; // @[MUL.scala 102:19]
  wire  m_1032_io_x3; // @[MUL.scala 102:19]
  wire  m_1032_io_s; // @[MUL.scala 102:19]
  wire  m_1032_io_cout; // @[MUL.scala 102:19]
  wire  m_1033_io_x1; // @[MUL.scala 102:19]
  wire  m_1033_io_x2; // @[MUL.scala 102:19]
  wire  m_1033_io_x3; // @[MUL.scala 102:19]
  wire  m_1033_io_s; // @[MUL.scala 102:19]
  wire  m_1033_io_cout; // @[MUL.scala 102:19]
  wire  m_1034_io_x1; // @[MUL.scala 102:19]
  wire  m_1034_io_x2; // @[MUL.scala 102:19]
  wire  m_1034_io_x3; // @[MUL.scala 102:19]
  wire  m_1034_io_s; // @[MUL.scala 102:19]
  wire  m_1034_io_cout; // @[MUL.scala 102:19]
  wire  m_1035_io_x1; // @[MUL.scala 102:19]
  wire  m_1035_io_x2; // @[MUL.scala 102:19]
  wire  m_1035_io_x3; // @[MUL.scala 102:19]
  wire  m_1035_io_s; // @[MUL.scala 102:19]
  wire  m_1035_io_cout; // @[MUL.scala 102:19]
  wire  m_1036_io_x1; // @[MUL.scala 102:19]
  wire  m_1036_io_x2; // @[MUL.scala 102:19]
  wire  m_1036_io_x3; // @[MUL.scala 102:19]
  wire  m_1036_io_s; // @[MUL.scala 102:19]
  wire  m_1036_io_cout; // @[MUL.scala 102:19]
  wire  m_1037_io_x1; // @[MUL.scala 102:19]
  wire  m_1037_io_x2; // @[MUL.scala 102:19]
  wire  m_1037_io_x3; // @[MUL.scala 102:19]
  wire  m_1037_io_s; // @[MUL.scala 102:19]
  wire  m_1037_io_cout; // @[MUL.scala 102:19]
  wire  m_1038_io_x1; // @[MUL.scala 102:19]
  wire  m_1038_io_x2; // @[MUL.scala 102:19]
  wire  m_1038_io_x3; // @[MUL.scala 102:19]
  wire  m_1038_io_s; // @[MUL.scala 102:19]
  wire  m_1038_io_cout; // @[MUL.scala 102:19]
  wire  m_1039_io_x1; // @[MUL.scala 102:19]
  wire  m_1039_io_x2; // @[MUL.scala 102:19]
  wire  m_1039_io_x3; // @[MUL.scala 102:19]
  wire  m_1039_io_s; // @[MUL.scala 102:19]
  wire  m_1039_io_cout; // @[MUL.scala 102:19]
  wire  m_1040_io_x1; // @[MUL.scala 102:19]
  wire  m_1040_io_x2; // @[MUL.scala 102:19]
  wire  m_1040_io_x3; // @[MUL.scala 102:19]
  wire  m_1040_io_s; // @[MUL.scala 102:19]
  wire  m_1040_io_cout; // @[MUL.scala 102:19]
  wire  m_1041_io_x1; // @[MUL.scala 102:19]
  wire  m_1041_io_x2; // @[MUL.scala 102:19]
  wire  m_1041_io_x3; // @[MUL.scala 102:19]
  wire  m_1041_io_s; // @[MUL.scala 102:19]
  wire  m_1041_io_cout; // @[MUL.scala 102:19]
  wire  m_1042_io_x1; // @[MUL.scala 102:19]
  wire  m_1042_io_x2; // @[MUL.scala 102:19]
  wire  m_1042_io_x3; // @[MUL.scala 102:19]
  wire  m_1042_io_s; // @[MUL.scala 102:19]
  wire  m_1042_io_cout; // @[MUL.scala 102:19]
  wire  m_1043_io_x1; // @[MUL.scala 102:19]
  wire  m_1043_io_x2; // @[MUL.scala 102:19]
  wire  m_1043_io_x3; // @[MUL.scala 102:19]
  wire  m_1043_io_s; // @[MUL.scala 102:19]
  wire  m_1043_io_cout; // @[MUL.scala 102:19]
  wire  m_1044_io_x1; // @[MUL.scala 102:19]
  wire  m_1044_io_x2; // @[MUL.scala 102:19]
  wire  m_1044_io_x3; // @[MUL.scala 102:19]
  wire  m_1044_io_s; // @[MUL.scala 102:19]
  wire  m_1044_io_cout; // @[MUL.scala 102:19]
  wire  m_1045_io_x1; // @[MUL.scala 102:19]
  wire  m_1045_io_x2; // @[MUL.scala 102:19]
  wire  m_1045_io_x3; // @[MUL.scala 102:19]
  wire  m_1045_io_s; // @[MUL.scala 102:19]
  wire  m_1045_io_cout; // @[MUL.scala 102:19]
  wire  m_1046_io_x1; // @[MUL.scala 102:19]
  wire  m_1046_io_x2; // @[MUL.scala 102:19]
  wire  m_1046_io_x3; // @[MUL.scala 102:19]
  wire  m_1046_io_s; // @[MUL.scala 102:19]
  wire  m_1046_io_cout; // @[MUL.scala 102:19]
  wire  m_1047_io_x1; // @[MUL.scala 102:19]
  wire  m_1047_io_x2; // @[MUL.scala 102:19]
  wire  m_1047_io_x3; // @[MUL.scala 102:19]
  wire  m_1047_io_s; // @[MUL.scala 102:19]
  wire  m_1047_io_cout; // @[MUL.scala 102:19]
  wire  m_1048_io_x1; // @[MUL.scala 102:19]
  wire  m_1048_io_x2; // @[MUL.scala 102:19]
  wire  m_1048_io_x3; // @[MUL.scala 102:19]
  wire  m_1048_io_s; // @[MUL.scala 102:19]
  wire  m_1048_io_cout; // @[MUL.scala 102:19]
  wire  m_1049_io_x1; // @[MUL.scala 102:19]
  wire  m_1049_io_x2; // @[MUL.scala 102:19]
  wire  m_1049_io_x3; // @[MUL.scala 102:19]
  wire  m_1049_io_s; // @[MUL.scala 102:19]
  wire  m_1049_io_cout; // @[MUL.scala 102:19]
  wire  m_1050_io_x1; // @[MUL.scala 102:19]
  wire  m_1050_io_x2; // @[MUL.scala 102:19]
  wire  m_1050_io_x3; // @[MUL.scala 102:19]
  wire  m_1050_io_s; // @[MUL.scala 102:19]
  wire  m_1050_io_cout; // @[MUL.scala 102:19]
  wire  m_1051_io_x1; // @[MUL.scala 102:19]
  wire  m_1051_io_x2; // @[MUL.scala 102:19]
  wire  m_1051_io_x3; // @[MUL.scala 102:19]
  wire  m_1051_io_s; // @[MUL.scala 102:19]
  wire  m_1051_io_cout; // @[MUL.scala 102:19]
  wire  m_1052_io_x1; // @[MUL.scala 102:19]
  wire  m_1052_io_x2; // @[MUL.scala 102:19]
  wire  m_1052_io_x3; // @[MUL.scala 102:19]
  wire  m_1052_io_s; // @[MUL.scala 102:19]
  wire  m_1052_io_cout; // @[MUL.scala 102:19]
  wire  m_1053_io_x1; // @[MUL.scala 102:19]
  wire  m_1053_io_x2; // @[MUL.scala 102:19]
  wire  m_1053_io_x3; // @[MUL.scala 102:19]
  wire  m_1053_io_s; // @[MUL.scala 102:19]
  wire  m_1053_io_cout; // @[MUL.scala 102:19]
  wire  m_1054_io_x1; // @[MUL.scala 102:19]
  wire  m_1054_io_x2; // @[MUL.scala 102:19]
  wire  m_1054_io_x3; // @[MUL.scala 102:19]
  wire  m_1054_io_s; // @[MUL.scala 102:19]
  wire  m_1054_io_cout; // @[MUL.scala 102:19]
  wire  m_1055_io_x1; // @[MUL.scala 102:19]
  wire  m_1055_io_x2; // @[MUL.scala 102:19]
  wire  m_1055_io_x3; // @[MUL.scala 102:19]
  wire  m_1055_io_s; // @[MUL.scala 102:19]
  wire  m_1055_io_cout; // @[MUL.scala 102:19]
  wire  m_1056_io_x1; // @[MUL.scala 102:19]
  wire  m_1056_io_x2; // @[MUL.scala 102:19]
  wire  m_1056_io_x3; // @[MUL.scala 102:19]
  wire  m_1056_io_s; // @[MUL.scala 102:19]
  wire  m_1056_io_cout; // @[MUL.scala 102:19]
  wire  m_1057_io_x1; // @[MUL.scala 102:19]
  wire  m_1057_io_x2; // @[MUL.scala 102:19]
  wire  m_1057_io_x3; // @[MUL.scala 102:19]
  wire  m_1057_io_s; // @[MUL.scala 102:19]
  wire  m_1057_io_cout; // @[MUL.scala 102:19]
  wire  m_1058_io_x1; // @[MUL.scala 102:19]
  wire  m_1058_io_x2; // @[MUL.scala 102:19]
  wire  m_1058_io_x3; // @[MUL.scala 102:19]
  wire  m_1058_io_s; // @[MUL.scala 102:19]
  wire  m_1058_io_cout; // @[MUL.scala 102:19]
  wire  m_1059_io_x1; // @[MUL.scala 102:19]
  wire  m_1059_io_x2; // @[MUL.scala 102:19]
  wire  m_1059_io_x3; // @[MUL.scala 102:19]
  wire  m_1059_io_s; // @[MUL.scala 102:19]
  wire  m_1059_io_cout; // @[MUL.scala 102:19]
  wire  m_1060_io_x1; // @[MUL.scala 102:19]
  wire  m_1060_io_x2; // @[MUL.scala 102:19]
  wire  m_1060_io_x3; // @[MUL.scala 102:19]
  wire  m_1060_io_s; // @[MUL.scala 102:19]
  wire  m_1060_io_cout; // @[MUL.scala 102:19]
  wire  m_1061_io_x1; // @[MUL.scala 102:19]
  wire  m_1061_io_x2; // @[MUL.scala 102:19]
  wire  m_1061_io_x3; // @[MUL.scala 102:19]
  wire  m_1061_io_s; // @[MUL.scala 102:19]
  wire  m_1061_io_cout; // @[MUL.scala 102:19]
  wire  m_1062_io_x1; // @[MUL.scala 102:19]
  wire  m_1062_io_x2; // @[MUL.scala 102:19]
  wire  m_1062_io_x3; // @[MUL.scala 102:19]
  wire  m_1062_io_s; // @[MUL.scala 102:19]
  wire  m_1062_io_cout; // @[MUL.scala 102:19]
  wire  m_1063_io_x1; // @[MUL.scala 102:19]
  wire  m_1063_io_x2; // @[MUL.scala 102:19]
  wire  m_1063_io_x3; // @[MUL.scala 102:19]
  wire  m_1063_io_s; // @[MUL.scala 102:19]
  wire  m_1063_io_cout; // @[MUL.scala 102:19]
  wire  m_1064_io_x1; // @[MUL.scala 102:19]
  wire  m_1064_io_x2; // @[MUL.scala 102:19]
  wire  m_1064_io_x3; // @[MUL.scala 102:19]
  wire  m_1064_io_s; // @[MUL.scala 102:19]
  wire  m_1064_io_cout; // @[MUL.scala 102:19]
  wire  m_1065_io_x1; // @[MUL.scala 102:19]
  wire  m_1065_io_x2; // @[MUL.scala 102:19]
  wire  m_1065_io_x3; // @[MUL.scala 102:19]
  wire  m_1065_io_s; // @[MUL.scala 102:19]
  wire  m_1065_io_cout; // @[MUL.scala 102:19]
  wire  m_1066_io_x1; // @[MUL.scala 102:19]
  wire  m_1066_io_x2; // @[MUL.scala 102:19]
  wire  m_1066_io_x3; // @[MUL.scala 102:19]
  wire  m_1066_io_s; // @[MUL.scala 102:19]
  wire  m_1066_io_cout; // @[MUL.scala 102:19]
  wire  m_1067_io_x1; // @[MUL.scala 102:19]
  wire  m_1067_io_x2; // @[MUL.scala 102:19]
  wire  m_1067_io_x3; // @[MUL.scala 102:19]
  wire  m_1067_io_s; // @[MUL.scala 102:19]
  wire  m_1067_io_cout; // @[MUL.scala 102:19]
  wire  m_1068_io_x1; // @[MUL.scala 102:19]
  wire  m_1068_io_x2; // @[MUL.scala 102:19]
  wire  m_1068_io_x3; // @[MUL.scala 102:19]
  wire  m_1068_io_s; // @[MUL.scala 102:19]
  wire  m_1068_io_cout; // @[MUL.scala 102:19]
  wire  m_1069_io_x1; // @[MUL.scala 102:19]
  wire  m_1069_io_x2; // @[MUL.scala 102:19]
  wire  m_1069_io_x3; // @[MUL.scala 102:19]
  wire  m_1069_io_s; // @[MUL.scala 102:19]
  wire  m_1069_io_cout; // @[MUL.scala 102:19]
  wire  m_1070_io_x1; // @[MUL.scala 102:19]
  wire  m_1070_io_x2; // @[MUL.scala 102:19]
  wire  m_1070_io_x3; // @[MUL.scala 102:19]
  wire  m_1070_io_s; // @[MUL.scala 102:19]
  wire  m_1070_io_cout; // @[MUL.scala 102:19]
  wire  m_1071_io_x1; // @[MUL.scala 102:19]
  wire  m_1071_io_x2; // @[MUL.scala 102:19]
  wire  m_1071_io_x3; // @[MUL.scala 102:19]
  wire  m_1071_io_s; // @[MUL.scala 102:19]
  wire  m_1071_io_cout; // @[MUL.scala 102:19]
  wire  m_1072_io_x1; // @[MUL.scala 102:19]
  wire  m_1072_io_x2; // @[MUL.scala 102:19]
  wire  m_1072_io_x3; // @[MUL.scala 102:19]
  wire  m_1072_io_s; // @[MUL.scala 102:19]
  wire  m_1072_io_cout; // @[MUL.scala 102:19]
  wire  m_1073_io_x1; // @[MUL.scala 102:19]
  wire  m_1073_io_x2; // @[MUL.scala 102:19]
  wire  m_1073_io_x3; // @[MUL.scala 102:19]
  wire  m_1073_io_s; // @[MUL.scala 102:19]
  wire  m_1073_io_cout; // @[MUL.scala 102:19]
  wire  m_1074_io_x1; // @[MUL.scala 102:19]
  wire  m_1074_io_x2; // @[MUL.scala 102:19]
  wire  m_1074_io_x3; // @[MUL.scala 102:19]
  wire  m_1074_io_s; // @[MUL.scala 102:19]
  wire  m_1074_io_cout; // @[MUL.scala 102:19]
  wire  m_1075_io_x1; // @[MUL.scala 102:19]
  wire  m_1075_io_x2; // @[MUL.scala 102:19]
  wire  m_1075_io_x3; // @[MUL.scala 102:19]
  wire  m_1075_io_s; // @[MUL.scala 102:19]
  wire  m_1075_io_cout; // @[MUL.scala 102:19]
  wire  m_1076_io_x1; // @[MUL.scala 102:19]
  wire  m_1076_io_x2; // @[MUL.scala 102:19]
  wire  m_1076_io_x3; // @[MUL.scala 102:19]
  wire  m_1076_io_s; // @[MUL.scala 102:19]
  wire  m_1076_io_cout; // @[MUL.scala 102:19]
  wire  m_1077_io_x1; // @[MUL.scala 102:19]
  wire  m_1077_io_x2; // @[MUL.scala 102:19]
  wire  m_1077_io_x3; // @[MUL.scala 102:19]
  wire  m_1077_io_s; // @[MUL.scala 102:19]
  wire  m_1077_io_cout; // @[MUL.scala 102:19]
  wire  m_1078_io_x1; // @[MUL.scala 102:19]
  wire  m_1078_io_x2; // @[MUL.scala 102:19]
  wire  m_1078_io_x3; // @[MUL.scala 102:19]
  wire  m_1078_io_s; // @[MUL.scala 102:19]
  wire  m_1078_io_cout; // @[MUL.scala 102:19]
  wire  m_1079_io_x1; // @[MUL.scala 102:19]
  wire  m_1079_io_x2; // @[MUL.scala 102:19]
  wire  m_1079_io_x3; // @[MUL.scala 102:19]
  wire  m_1079_io_s; // @[MUL.scala 102:19]
  wire  m_1079_io_cout; // @[MUL.scala 102:19]
  wire  m_1080_io_x1; // @[MUL.scala 102:19]
  wire  m_1080_io_x2; // @[MUL.scala 102:19]
  wire  m_1080_io_x3; // @[MUL.scala 102:19]
  wire  m_1080_io_s; // @[MUL.scala 102:19]
  wire  m_1080_io_cout; // @[MUL.scala 102:19]
  wire  m_1081_io_x1; // @[MUL.scala 102:19]
  wire  m_1081_io_x2; // @[MUL.scala 102:19]
  wire  m_1081_io_x3; // @[MUL.scala 102:19]
  wire  m_1081_io_s; // @[MUL.scala 102:19]
  wire  m_1081_io_cout; // @[MUL.scala 102:19]
  wire  m_1082_io_x1; // @[MUL.scala 102:19]
  wire  m_1082_io_x2; // @[MUL.scala 102:19]
  wire  m_1082_io_x3; // @[MUL.scala 102:19]
  wire  m_1082_io_s; // @[MUL.scala 102:19]
  wire  m_1082_io_cout; // @[MUL.scala 102:19]
  wire  m_1083_io_x1; // @[MUL.scala 102:19]
  wire  m_1083_io_x2; // @[MUL.scala 102:19]
  wire  m_1083_io_x3; // @[MUL.scala 102:19]
  wire  m_1083_io_s; // @[MUL.scala 102:19]
  wire  m_1083_io_cout; // @[MUL.scala 102:19]
  wire  m_1084_io_x1; // @[MUL.scala 102:19]
  wire  m_1084_io_x2; // @[MUL.scala 102:19]
  wire  m_1084_io_x3; // @[MUL.scala 102:19]
  wire  m_1084_io_s; // @[MUL.scala 102:19]
  wire  m_1084_io_cout; // @[MUL.scala 102:19]
  wire  m_1085_io_x1; // @[MUL.scala 102:19]
  wire  m_1085_io_x2; // @[MUL.scala 102:19]
  wire  m_1085_io_x3; // @[MUL.scala 102:19]
  wire  m_1085_io_s; // @[MUL.scala 102:19]
  wire  m_1085_io_cout; // @[MUL.scala 102:19]
  wire  m_1086_io_x1; // @[MUL.scala 102:19]
  wire  m_1086_io_x2; // @[MUL.scala 102:19]
  wire  m_1086_io_x3; // @[MUL.scala 102:19]
  wire  m_1086_io_s; // @[MUL.scala 102:19]
  wire  m_1086_io_cout; // @[MUL.scala 102:19]
  wire  m_1087_io_x1; // @[MUL.scala 102:19]
  wire  m_1087_io_x2; // @[MUL.scala 102:19]
  wire  m_1087_io_x3; // @[MUL.scala 102:19]
  wire  m_1087_io_s; // @[MUL.scala 102:19]
  wire  m_1087_io_cout; // @[MUL.scala 102:19]
  wire  m_1088_io_x1; // @[MUL.scala 102:19]
  wire  m_1088_io_x2; // @[MUL.scala 102:19]
  wire  m_1088_io_x3; // @[MUL.scala 102:19]
  wire  m_1088_io_s; // @[MUL.scala 102:19]
  wire  m_1088_io_cout; // @[MUL.scala 102:19]
  wire  m_1089_io_x1; // @[MUL.scala 102:19]
  wire  m_1089_io_x2; // @[MUL.scala 102:19]
  wire  m_1089_io_x3; // @[MUL.scala 102:19]
  wire  m_1089_io_s; // @[MUL.scala 102:19]
  wire  m_1089_io_cout; // @[MUL.scala 102:19]
  wire  m_1090_io_x1; // @[MUL.scala 102:19]
  wire  m_1090_io_x2; // @[MUL.scala 102:19]
  wire  m_1090_io_x3; // @[MUL.scala 102:19]
  wire  m_1090_io_s; // @[MUL.scala 102:19]
  wire  m_1090_io_cout; // @[MUL.scala 102:19]
  wire  m_1091_io_x1; // @[MUL.scala 102:19]
  wire  m_1091_io_x2; // @[MUL.scala 102:19]
  wire  m_1091_io_x3; // @[MUL.scala 102:19]
  wire  m_1091_io_s; // @[MUL.scala 102:19]
  wire  m_1091_io_cout; // @[MUL.scala 102:19]
  wire  m_1092_io_x1; // @[MUL.scala 102:19]
  wire  m_1092_io_x2; // @[MUL.scala 102:19]
  wire  m_1092_io_x3; // @[MUL.scala 102:19]
  wire  m_1092_io_s; // @[MUL.scala 102:19]
  wire  m_1092_io_cout; // @[MUL.scala 102:19]
  wire  m_1093_io_x1; // @[MUL.scala 102:19]
  wire  m_1093_io_x2; // @[MUL.scala 102:19]
  wire  m_1093_io_x3; // @[MUL.scala 102:19]
  wire  m_1093_io_s; // @[MUL.scala 102:19]
  wire  m_1093_io_cout; // @[MUL.scala 102:19]
  wire  m_1094_io_x1; // @[MUL.scala 102:19]
  wire  m_1094_io_x2; // @[MUL.scala 102:19]
  wire  m_1094_io_x3; // @[MUL.scala 102:19]
  wire  m_1094_io_s; // @[MUL.scala 102:19]
  wire  m_1094_io_cout; // @[MUL.scala 102:19]
  wire  m_1095_io_x1; // @[MUL.scala 102:19]
  wire  m_1095_io_x2; // @[MUL.scala 102:19]
  wire  m_1095_io_x3; // @[MUL.scala 102:19]
  wire  m_1095_io_s; // @[MUL.scala 102:19]
  wire  m_1095_io_cout; // @[MUL.scala 102:19]
  wire  m_1096_io_x1; // @[MUL.scala 102:19]
  wire  m_1096_io_x2; // @[MUL.scala 102:19]
  wire  m_1096_io_x3; // @[MUL.scala 102:19]
  wire  m_1096_io_s; // @[MUL.scala 102:19]
  wire  m_1096_io_cout; // @[MUL.scala 102:19]
  wire  m_1097_io_x1; // @[MUL.scala 102:19]
  wire  m_1097_io_x2; // @[MUL.scala 102:19]
  wire  m_1097_io_x3; // @[MUL.scala 102:19]
  wire  m_1097_io_s; // @[MUL.scala 102:19]
  wire  m_1097_io_cout; // @[MUL.scala 102:19]
  wire  m_1098_io_x1; // @[MUL.scala 102:19]
  wire  m_1098_io_x2; // @[MUL.scala 102:19]
  wire  m_1098_io_x3; // @[MUL.scala 102:19]
  wire  m_1098_io_s; // @[MUL.scala 102:19]
  wire  m_1098_io_cout; // @[MUL.scala 102:19]
  wire  m_1099_io_x1; // @[MUL.scala 102:19]
  wire  m_1099_io_x2; // @[MUL.scala 102:19]
  wire  m_1099_io_x3; // @[MUL.scala 102:19]
  wire  m_1099_io_s; // @[MUL.scala 102:19]
  wire  m_1099_io_cout; // @[MUL.scala 102:19]
  wire  m_1100_io_x1; // @[MUL.scala 102:19]
  wire  m_1100_io_x2; // @[MUL.scala 102:19]
  wire  m_1100_io_x3; // @[MUL.scala 102:19]
  wire  m_1100_io_s; // @[MUL.scala 102:19]
  wire  m_1100_io_cout; // @[MUL.scala 102:19]
  wire  m_1101_io_x1; // @[MUL.scala 102:19]
  wire  m_1101_io_x2; // @[MUL.scala 102:19]
  wire  m_1101_io_x3; // @[MUL.scala 102:19]
  wire  m_1101_io_s; // @[MUL.scala 102:19]
  wire  m_1101_io_cout; // @[MUL.scala 102:19]
  wire  m_1102_io_x1; // @[MUL.scala 102:19]
  wire  m_1102_io_x2; // @[MUL.scala 102:19]
  wire  m_1102_io_x3; // @[MUL.scala 102:19]
  wire  m_1102_io_s; // @[MUL.scala 102:19]
  wire  m_1102_io_cout; // @[MUL.scala 102:19]
  wire  m_1103_io_x1; // @[MUL.scala 102:19]
  wire  m_1103_io_x2; // @[MUL.scala 102:19]
  wire  m_1103_io_x3; // @[MUL.scala 102:19]
  wire  m_1103_io_s; // @[MUL.scala 102:19]
  wire  m_1103_io_cout; // @[MUL.scala 102:19]
  wire  m_1104_io_x1; // @[MUL.scala 102:19]
  wire  m_1104_io_x2; // @[MUL.scala 102:19]
  wire  m_1104_io_x3; // @[MUL.scala 102:19]
  wire  m_1104_io_s; // @[MUL.scala 102:19]
  wire  m_1104_io_cout; // @[MUL.scala 102:19]
  wire  m_1105_io_x1; // @[MUL.scala 102:19]
  wire  m_1105_io_x2; // @[MUL.scala 102:19]
  wire  m_1105_io_x3; // @[MUL.scala 102:19]
  wire  m_1105_io_s; // @[MUL.scala 102:19]
  wire  m_1105_io_cout; // @[MUL.scala 102:19]
  wire  m_1106_io_x1; // @[MUL.scala 102:19]
  wire  m_1106_io_x2; // @[MUL.scala 102:19]
  wire  m_1106_io_x3; // @[MUL.scala 102:19]
  wire  m_1106_io_s; // @[MUL.scala 102:19]
  wire  m_1106_io_cout; // @[MUL.scala 102:19]
  wire  m_1107_io_x1; // @[MUL.scala 102:19]
  wire  m_1107_io_x2; // @[MUL.scala 102:19]
  wire  m_1107_io_x3; // @[MUL.scala 102:19]
  wire  m_1107_io_s; // @[MUL.scala 102:19]
  wire  m_1107_io_cout; // @[MUL.scala 102:19]
  wire  m_1108_io_x1; // @[MUL.scala 102:19]
  wire  m_1108_io_x2; // @[MUL.scala 102:19]
  wire  m_1108_io_x3; // @[MUL.scala 102:19]
  wire  m_1108_io_s; // @[MUL.scala 102:19]
  wire  m_1108_io_cout; // @[MUL.scala 102:19]
  wire  m_1109_io_x1; // @[MUL.scala 102:19]
  wire  m_1109_io_x2; // @[MUL.scala 102:19]
  wire  m_1109_io_x3; // @[MUL.scala 102:19]
  wire  m_1109_io_s; // @[MUL.scala 102:19]
  wire  m_1109_io_cout; // @[MUL.scala 102:19]
  wire  m_1110_io_x1; // @[MUL.scala 102:19]
  wire  m_1110_io_x2; // @[MUL.scala 102:19]
  wire  m_1110_io_x3; // @[MUL.scala 102:19]
  wire  m_1110_io_s; // @[MUL.scala 102:19]
  wire  m_1110_io_cout; // @[MUL.scala 102:19]
  wire  m_1111_io_x1; // @[MUL.scala 102:19]
  wire  m_1111_io_x2; // @[MUL.scala 102:19]
  wire  m_1111_io_x3; // @[MUL.scala 102:19]
  wire  m_1111_io_s; // @[MUL.scala 102:19]
  wire  m_1111_io_cout; // @[MUL.scala 102:19]
  wire  m_1112_io_x1; // @[MUL.scala 102:19]
  wire  m_1112_io_x2; // @[MUL.scala 102:19]
  wire  m_1112_io_x3; // @[MUL.scala 102:19]
  wire  m_1112_io_s; // @[MUL.scala 102:19]
  wire  m_1112_io_cout; // @[MUL.scala 102:19]
  wire  m_1113_io_x1; // @[MUL.scala 102:19]
  wire  m_1113_io_x2; // @[MUL.scala 102:19]
  wire  m_1113_io_x3; // @[MUL.scala 102:19]
  wire  m_1113_io_s; // @[MUL.scala 102:19]
  wire  m_1113_io_cout; // @[MUL.scala 102:19]
  wire  m_1114_io_x1; // @[MUL.scala 102:19]
  wire  m_1114_io_x2; // @[MUL.scala 102:19]
  wire  m_1114_io_x3; // @[MUL.scala 102:19]
  wire  m_1114_io_s; // @[MUL.scala 102:19]
  wire  m_1114_io_cout; // @[MUL.scala 102:19]
  wire  m_1115_io_x1; // @[MUL.scala 102:19]
  wire  m_1115_io_x2; // @[MUL.scala 102:19]
  wire  m_1115_io_x3; // @[MUL.scala 102:19]
  wire  m_1115_io_s; // @[MUL.scala 102:19]
  wire  m_1115_io_cout; // @[MUL.scala 102:19]
  wire  m_1116_io_x1; // @[MUL.scala 102:19]
  wire  m_1116_io_x2; // @[MUL.scala 102:19]
  wire  m_1116_io_x3; // @[MUL.scala 102:19]
  wire  m_1116_io_s; // @[MUL.scala 102:19]
  wire  m_1116_io_cout; // @[MUL.scala 102:19]
  wire  m_1117_io_in_0; // @[MUL.scala 124:19]
  wire  m_1117_io_in_1; // @[MUL.scala 124:19]
  wire  m_1117_io_out_0; // @[MUL.scala 124:19]
  wire  m_1117_io_out_1; // @[MUL.scala 124:19]
  wire  m_1118_io_x1; // @[MUL.scala 102:19]
  wire  m_1118_io_x2; // @[MUL.scala 102:19]
  wire  m_1118_io_x3; // @[MUL.scala 102:19]
  wire  m_1118_io_s; // @[MUL.scala 102:19]
  wire  m_1118_io_cout; // @[MUL.scala 102:19]
  wire  m_1119_io_x1; // @[MUL.scala 102:19]
  wire  m_1119_io_x2; // @[MUL.scala 102:19]
  wire  m_1119_io_x3; // @[MUL.scala 102:19]
  wire  m_1119_io_s; // @[MUL.scala 102:19]
  wire  m_1119_io_cout; // @[MUL.scala 102:19]
  wire  m_1120_io_x1; // @[MUL.scala 102:19]
  wire  m_1120_io_x2; // @[MUL.scala 102:19]
  wire  m_1120_io_x3; // @[MUL.scala 102:19]
  wire  m_1120_io_s; // @[MUL.scala 102:19]
  wire  m_1120_io_cout; // @[MUL.scala 102:19]
  wire  m_1121_io_x1; // @[MUL.scala 102:19]
  wire  m_1121_io_x2; // @[MUL.scala 102:19]
  wire  m_1121_io_x3; // @[MUL.scala 102:19]
  wire  m_1121_io_s; // @[MUL.scala 102:19]
  wire  m_1121_io_cout; // @[MUL.scala 102:19]
  wire  m_1122_io_x1; // @[MUL.scala 102:19]
  wire  m_1122_io_x2; // @[MUL.scala 102:19]
  wire  m_1122_io_x3; // @[MUL.scala 102:19]
  wire  m_1122_io_s; // @[MUL.scala 102:19]
  wire  m_1122_io_cout; // @[MUL.scala 102:19]
  wire  m_1123_io_x1; // @[MUL.scala 102:19]
  wire  m_1123_io_x2; // @[MUL.scala 102:19]
  wire  m_1123_io_x3; // @[MUL.scala 102:19]
  wire  m_1123_io_s; // @[MUL.scala 102:19]
  wire  m_1123_io_cout; // @[MUL.scala 102:19]
  wire  m_1124_io_in_0; // @[MUL.scala 124:19]
  wire  m_1124_io_in_1; // @[MUL.scala 124:19]
  wire  m_1124_io_out_0; // @[MUL.scala 124:19]
  wire  m_1124_io_out_1; // @[MUL.scala 124:19]
  wire  m_1125_io_x1; // @[MUL.scala 102:19]
  wire  m_1125_io_x2; // @[MUL.scala 102:19]
  wire  m_1125_io_x3; // @[MUL.scala 102:19]
  wire  m_1125_io_s; // @[MUL.scala 102:19]
  wire  m_1125_io_cout; // @[MUL.scala 102:19]
  wire  m_1126_io_x1; // @[MUL.scala 102:19]
  wire  m_1126_io_x2; // @[MUL.scala 102:19]
  wire  m_1126_io_x3; // @[MUL.scala 102:19]
  wire  m_1126_io_s; // @[MUL.scala 102:19]
  wire  m_1126_io_cout; // @[MUL.scala 102:19]
  wire  m_1127_io_x1; // @[MUL.scala 102:19]
  wire  m_1127_io_x2; // @[MUL.scala 102:19]
  wire  m_1127_io_x3; // @[MUL.scala 102:19]
  wire  m_1127_io_s; // @[MUL.scala 102:19]
  wire  m_1127_io_cout; // @[MUL.scala 102:19]
  wire  m_1128_io_x1; // @[MUL.scala 102:19]
  wire  m_1128_io_x2; // @[MUL.scala 102:19]
  wire  m_1128_io_x3; // @[MUL.scala 102:19]
  wire  m_1128_io_s; // @[MUL.scala 102:19]
  wire  m_1128_io_cout; // @[MUL.scala 102:19]
  wire  m_1129_io_x1; // @[MUL.scala 102:19]
  wire  m_1129_io_x2; // @[MUL.scala 102:19]
  wire  m_1129_io_x3; // @[MUL.scala 102:19]
  wire  m_1129_io_s; // @[MUL.scala 102:19]
  wire  m_1129_io_cout; // @[MUL.scala 102:19]
  wire  m_1130_io_x1; // @[MUL.scala 102:19]
  wire  m_1130_io_x2; // @[MUL.scala 102:19]
  wire  m_1130_io_x3; // @[MUL.scala 102:19]
  wire  m_1130_io_s; // @[MUL.scala 102:19]
  wire  m_1130_io_cout; // @[MUL.scala 102:19]
  wire  m_1131_io_in_0; // @[MUL.scala 124:19]
  wire  m_1131_io_in_1; // @[MUL.scala 124:19]
  wire  m_1131_io_out_0; // @[MUL.scala 124:19]
  wire  m_1131_io_out_1; // @[MUL.scala 124:19]
  wire  m_1132_io_x1; // @[MUL.scala 102:19]
  wire  m_1132_io_x2; // @[MUL.scala 102:19]
  wire  m_1132_io_x3; // @[MUL.scala 102:19]
  wire  m_1132_io_s; // @[MUL.scala 102:19]
  wire  m_1132_io_cout; // @[MUL.scala 102:19]
  wire  m_1133_io_x1; // @[MUL.scala 102:19]
  wire  m_1133_io_x2; // @[MUL.scala 102:19]
  wire  m_1133_io_x3; // @[MUL.scala 102:19]
  wire  m_1133_io_s; // @[MUL.scala 102:19]
  wire  m_1133_io_cout; // @[MUL.scala 102:19]
  wire  m_1134_io_x1; // @[MUL.scala 102:19]
  wire  m_1134_io_x2; // @[MUL.scala 102:19]
  wire  m_1134_io_x3; // @[MUL.scala 102:19]
  wire  m_1134_io_s; // @[MUL.scala 102:19]
  wire  m_1134_io_cout; // @[MUL.scala 102:19]
  wire  m_1135_io_x1; // @[MUL.scala 102:19]
  wire  m_1135_io_x2; // @[MUL.scala 102:19]
  wire  m_1135_io_x3; // @[MUL.scala 102:19]
  wire  m_1135_io_s; // @[MUL.scala 102:19]
  wire  m_1135_io_cout; // @[MUL.scala 102:19]
  wire  m_1136_io_x1; // @[MUL.scala 102:19]
  wire  m_1136_io_x2; // @[MUL.scala 102:19]
  wire  m_1136_io_x3; // @[MUL.scala 102:19]
  wire  m_1136_io_s; // @[MUL.scala 102:19]
  wire  m_1136_io_cout; // @[MUL.scala 102:19]
  wire  m_1137_io_x1; // @[MUL.scala 102:19]
  wire  m_1137_io_x2; // @[MUL.scala 102:19]
  wire  m_1137_io_x3; // @[MUL.scala 102:19]
  wire  m_1137_io_s; // @[MUL.scala 102:19]
  wire  m_1137_io_cout; // @[MUL.scala 102:19]
  wire  m_1138_io_in_0; // @[MUL.scala 124:19]
  wire  m_1138_io_in_1; // @[MUL.scala 124:19]
  wire  m_1138_io_out_0; // @[MUL.scala 124:19]
  wire  m_1138_io_out_1; // @[MUL.scala 124:19]
  wire  m_1139_io_x1; // @[MUL.scala 102:19]
  wire  m_1139_io_x2; // @[MUL.scala 102:19]
  wire  m_1139_io_x3; // @[MUL.scala 102:19]
  wire  m_1139_io_s; // @[MUL.scala 102:19]
  wire  m_1139_io_cout; // @[MUL.scala 102:19]
  wire  m_1140_io_x1; // @[MUL.scala 102:19]
  wire  m_1140_io_x2; // @[MUL.scala 102:19]
  wire  m_1140_io_x3; // @[MUL.scala 102:19]
  wire  m_1140_io_s; // @[MUL.scala 102:19]
  wire  m_1140_io_cout; // @[MUL.scala 102:19]
  wire  m_1141_io_x1; // @[MUL.scala 102:19]
  wire  m_1141_io_x2; // @[MUL.scala 102:19]
  wire  m_1141_io_x3; // @[MUL.scala 102:19]
  wire  m_1141_io_s; // @[MUL.scala 102:19]
  wire  m_1141_io_cout; // @[MUL.scala 102:19]
  wire  m_1142_io_x1; // @[MUL.scala 102:19]
  wire  m_1142_io_x2; // @[MUL.scala 102:19]
  wire  m_1142_io_x3; // @[MUL.scala 102:19]
  wire  m_1142_io_s; // @[MUL.scala 102:19]
  wire  m_1142_io_cout; // @[MUL.scala 102:19]
  wire  m_1143_io_x1; // @[MUL.scala 102:19]
  wire  m_1143_io_x2; // @[MUL.scala 102:19]
  wire  m_1143_io_x3; // @[MUL.scala 102:19]
  wire  m_1143_io_s; // @[MUL.scala 102:19]
  wire  m_1143_io_cout; // @[MUL.scala 102:19]
  wire  m_1144_io_x1; // @[MUL.scala 102:19]
  wire  m_1144_io_x2; // @[MUL.scala 102:19]
  wire  m_1144_io_x3; // @[MUL.scala 102:19]
  wire  m_1144_io_s; // @[MUL.scala 102:19]
  wire  m_1144_io_cout; // @[MUL.scala 102:19]
  wire  m_1145_io_in_0; // @[MUL.scala 124:19]
  wire  m_1145_io_in_1; // @[MUL.scala 124:19]
  wire  m_1145_io_out_0; // @[MUL.scala 124:19]
  wire  m_1145_io_out_1; // @[MUL.scala 124:19]
  wire  m_1146_io_x1; // @[MUL.scala 102:19]
  wire  m_1146_io_x2; // @[MUL.scala 102:19]
  wire  m_1146_io_x3; // @[MUL.scala 102:19]
  wire  m_1146_io_s; // @[MUL.scala 102:19]
  wire  m_1146_io_cout; // @[MUL.scala 102:19]
  wire  m_1147_io_x1; // @[MUL.scala 102:19]
  wire  m_1147_io_x2; // @[MUL.scala 102:19]
  wire  m_1147_io_x3; // @[MUL.scala 102:19]
  wire  m_1147_io_s; // @[MUL.scala 102:19]
  wire  m_1147_io_cout; // @[MUL.scala 102:19]
  wire  m_1148_io_x1; // @[MUL.scala 102:19]
  wire  m_1148_io_x2; // @[MUL.scala 102:19]
  wire  m_1148_io_x3; // @[MUL.scala 102:19]
  wire  m_1148_io_s; // @[MUL.scala 102:19]
  wire  m_1148_io_cout; // @[MUL.scala 102:19]
  wire  m_1149_io_x1; // @[MUL.scala 102:19]
  wire  m_1149_io_x2; // @[MUL.scala 102:19]
  wire  m_1149_io_x3; // @[MUL.scala 102:19]
  wire  m_1149_io_s; // @[MUL.scala 102:19]
  wire  m_1149_io_cout; // @[MUL.scala 102:19]
  wire  m_1150_io_x1; // @[MUL.scala 102:19]
  wire  m_1150_io_x2; // @[MUL.scala 102:19]
  wire  m_1150_io_x3; // @[MUL.scala 102:19]
  wire  m_1150_io_s; // @[MUL.scala 102:19]
  wire  m_1150_io_cout; // @[MUL.scala 102:19]
  wire  m_1151_io_x1; // @[MUL.scala 102:19]
  wire  m_1151_io_x2; // @[MUL.scala 102:19]
  wire  m_1151_io_x3; // @[MUL.scala 102:19]
  wire  m_1151_io_s; // @[MUL.scala 102:19]
  wire  m_1151_io_cout; // @[MUL.scala 102:19]
  wire  m_1152_io_x1; // @[MUL.scala 102:19]
  wire  m_1152_io_x2; // @[MUL.scala 102:19]
  wire  m_1152_io_x3; // @[MUL.scala 102:19]
  wire  m_1152_io_s; // @[MUL.scala 102:19]
  wire  m_1152_io_cout; // @[MUL.scala 102:19]
  wire  m_1153_io_x1; // @[MUL.scala 102:19]
  wire  m_1153_io_x2; // @[MUL.scala 102:19]
  wire  m_1153_io_x3; // @[MUL.scala 102:19]
  wire  m_1153_io_s; // @[MUL.scala 102:19]
  wire  m_1153_io_cout; // @[MUL.scala 102:19]
  wire  m_1154_io_x1; // @[MUL.scala 102:19]
  wire  m_1154_io_x2; // @[MUL.scala 102:19]
  wire  m_1154_io_x3; // @[MUL.scala 102:19]
  wire  m_1154_io_s; // @[MUL.scala 102:19]
  wire  m_1154_io_cout; // @[MUL.scala 102:19]
  wire  m_1155_io_x1; // @[MUL.scala 102:19]
  wire  m_1155_io_x2; // @[MUL.scala 102:19]
  wire  m_1155_io_x3; // @[MUL.scala 102:19]
  wire  m_1155_io_s; // @[MUL.scala 102:19]
  wire  m_1155_io_cout; // @[MUL.scala 102:19]
  wire  m_1156_io_x1; // @[MUL.scala 102:19]
  wire  m_1156_io_x2; // @[MUL.scala 102:19]
  wire  m_1156_io_x3; // @[MUL.scala 102:19]
  wire  m_1156_io_s; // @[MUL.scala 102:19]
  wire  m_1156_io_cout; // @[MUL.scala 102:19]
  wire  m_1157_io_x1; // @[MUL.scala 102:19]
  wire  m_1157_io_x2; // @[MUL.scala 102:19]
  wire  m_1157_io_x3; // @[MUL.scala 102:19]
  wire  m_1157_io_s; // @[MUL.scala 102:19]
  wire  m_1157_io_cout; // @[MUL.scala 102:19]
  wire  m_1158_io_x1; // @[MUL.scala 102:19]
  wire  m_1158_io_x2; // @[MUL.scala 102:19]
  wire  m_1158_io_x3; // @[MUL.scala 102:19]
  wire  m_1158_io_s; // @[MUL.scala 102:19]
  wire  m_1158_io_cout; // @[MUL.scala 102:19]
  wire  m_1159_io_x1; // @[MUL.scala 102:19]
  wire  m_1159_io_x2; // @[MUL.scala 102:19]
  wire  m_1159_io_x3; // @[MUL.scala 102:19]
  wire  m_1159_io_s; // @[MUL.scala 102:19]
  wire  m_1159_io_cout; // @[MUL.scala 102:19]
  wire  m_1160_io_x1; // @[MUL.scala 102:19]
  wire  m_1160_io_x2; // @[MUL.scala 102:19]
  wire  m_1160_io_x3; // @[MUL.scala 102:19]
  wire  m_1160_io_s; // @[MUL.scala 102:19]
  wire  m_1160_io_cout; // @[MUL.scala 102:19]
  wire  m_1161_io_x1; // @[MUL.scala 102:19]
  wire  m_1161_io_x2; // @[MUL.scala 102:19]
  wire  m_1161_io_x3; // @[MUL.scala 102:19]
  wire  m_1161_io_s; // @[MUL.scala 102:19]
  wire  m_1161_io_cout; // @[MUL.scala 102:19]
  wire  m_1162_io_x1; // @[MUL.scala 102:19]
  wire  m_1162_io_x2; // @[MUL.scala 102:19]
  wire  m_1162_io_x3; // @[MUL.scala 102:19]
  wire  m_1162_io_s; // @[MUL.scala 102:19]
  wire  m_1162_io_cout; // @[MUL.scala 102:19]
  wire  m_1163_io_x1; // @[MUL.scala 102:19]
  wire  m_1163_io_x2; // @[MUL.scala 102:19]
  wire  m_1163_io_x3; // @[MUL.scala 102:19]
  wire  m_1163_io_s; // @[MUL.scala 102:19]
  wire  m_1163_io_cout; // @[MUL.scala 102:19]
  wire  m_1164_io_x1; // @[MUL.scala 102:19]
  wire  m_1164_io_x2; // @[MUL.scala 102:19]
  wire  m_1164_io_x3; // @[MUL.scala 102:19]
  wire  m_1164_io_s; // @[MUL.scala 102:19]
  wire  m_1164_io_cout; // @[MUL.scala 102:19]
  wire  m_1165_io_x1; // @[MUL.scala 102:19]
  wire  m_1165_io_x2; // @[MUL.scala 102:19]
  wire  m_1165_io_x3; // @[MUL.scala 102:19]
  wire  m_1165_io_s; // @[MUL.scala 102:19]
  wire  m_1165_io_cout; // @[MUL.scala 102:19]
  wire  m_1166_io_x1; // @[MUL.scala 102:19]
  wire  m_1166_io_x2; // @[MUL.scala 102:19]
  wire  m_1166_io_x3; // @[MUL.scala 102:19]
  wire  m_1166_io_s; // @[MUL.scala 102:19]
  wire  m_1166_io_cout; // @[MUL.scala 102:19]
  wire  m_1167_io_x1; // @[MUL.scala 102:19]
  wire  m_1167_io_x2; // @[MUL.scala 102:19]
  wire  m_1167_io_x3; // @[MUL.scala 102:19]
  wire  m_1167_io_s; // @[MUL.scala 102:19]
  wire  m_1167_io_cout; // @[MUL.scala 102:19]
  wire  m_1168_io_x1; // @[MUL.scala 102:19]
  wire  m_1168_io_x2; // @[MUL.scala 102:19]
  wire  m_1168_io_x3; // @[MUL.scala 102:19]
  wire  m_1168_io_s; // @[MUL.scala 102:19]
  wire  m_1168_io_cout; // @[MUL.scala 102:19]
  wire  m_1169_io_x1; // @[MUL.scala 102:19]
  wire  m_1169_io_x2; // @[MUL.scala 102:19]
  wire  m_1169_io_x3; // @[MUL.scala 102:19]
  wire  m_1169_io_s; // @[MUL.scala 102:19]
  wire  m_1169_io_cout; // @[MUL.scala 102:19]
  wire  m_1170_io_x1; // @[MUL.scala 102:19]
  wire  m_1170_io_x2; // @[MUL.scala 102:19]
  wire  m_1170_io_x3; // @[MUL.scala 102:19]
  wire  m_1170_io_s; // @[MUL.scala 102:19]
  wire  m_1170_io_cout; // @[MUL.scala 102:19]
  wire  m_1171_io_x1; // @[MUL.scala 102:19]
  wire  m_1171_io_x2; // @[MUL.scala 102:19]
  wire  m_1171_io_x3; // @[MUL.scala 102:19]
  wire  m_1171_io_s; // @[MUL.scala 102:19]
  wire  m_1171_io_cout; // @[MUL.scala 102:19]
  wire  m_1172_io_x1; // @[MUL.scala 102:19]
  wire  m_1172_io_x2; // @[MUL.scala 102:19]
  wire  m_1172_io_x3; // @[MUL.scala 102:19]
  wire  m_1172_io_s; // @[MUL.scala 102:19]
  wire  m_1172_io_cout; // @[MUL.scala 102:19]
  wire  m_1173_io_x1; // @[MUL.scala 102:19]
  wire  m_1173_io_x2; // @[MUL.scala 102:19]
  wire  m_1173_io_x3; // @[MUL.scala 102:19]
  wire  m_1173_io_s; // @[MUL.scala 102:19]
  wire  m_1173_io_cout; // @[MUL.scala 102:19]
  wire  m_1174_io_x1; // @[MUL.scala 102:19]
  wire  m_1174_io_x2; // @[MUL.scala 102:19]
  wire  m_1174_io_x3; // @[MUL.scala 102:19]
  wire  m_1174_io_s; // @[MUL.scala 102:19]
  wire  m_1174_io_cout; // @[MUL.scala 102:19]
  wire  m_1175_io_x1; // @[MUL.scala 102:19]
  wire  m_1175_io_x2; // @[MUL.scala 102:19]
  wire  m_1175_io_x3; // @[MUL.scala 102:19]
  wire  m_1175_io_s; // @[MUL.scala 102:19]
  wire  m_1175_io_cout; // @[MUL.scala 102:19]
  wire  m_1176_io_x1; // @[MUL.scala 102:19]
  wire  m_1176_io_x2; // @[MUL.scala 102:19]
  wire  m_1176_io_x3; // @[MUL.scala 102:19]
  wire  m_1176_io_s; // @[MUL.scala 102:19]
  wire  m_1176_io_cout; // @[MUL.scala 102:19]
  wire  m_1177_io_x1; // @[MUL.scala 102:19]
  wire  m_1177_io_x2; // @[MUL.scala 102:19]
  wire  m_1177_io_x3; // @[MUL.scala 102:19]
  wire  m_1177_io_s; // @[MUL.scala 102:19]
  wire  m_1177_io_cout; // @[MUL.scala 102:19]
  wire  m_1178_io_x1; // @[MUL.scala 102:19]
  wire  m_1178_io_x2; // @[MUL.scala 102:19]
  wire  m_1178_io_x3; // @[MUL.scala 102:19]
  wire  m_1178_io_s; // @[MUL.scala 102:19]
  wire  m_1178_io_cout; // @[MUL.scala 102:19]
  wire  m_1179_io_x1; // @[MUL.scala 102:19]
  wire  m_1179_io_x2; // @[MUL.scala 102:19]
  wire  m_1179_io_x3; // @[MUL.scala 102:19]
  wire  m_1179_io_s; // @[MUL.scala 102:19]
  wire  m_1179_io_cout; // @[MUL.scala 102:19]
  wire  m_1180_io_x1; // @[MUL.scala 102:19]
  wire  m_1180_io_x2; // @[MUL.scala 102:19]
  wire  m_1180_io_x3; // @[MUL.scala 102:19]
  wire  m_1180_io_s; // @[MUL.scala 102:19]
  wire  m_1180_io_cout; // @[MUL.scala 102:19]
  wire  m_1181_io_x1; // @[MUL.scala 102:19]
  wire  m_1181_io_x2; // @[MUL.scala 102:19]
  wire  m_1181_io_x3; // @[MUL.scala 102:19]
  wire  m_1181_io_s; // @[MUL.scala 102:19]
  wire  m_1181_io_cout; // @[MUL.scala 102:19]
  wire  m_1182_io_x1; // @[MUL.scala 102:19]
  wire  m_1182_io_x2; // @[MUL.scala 102:19]
  wire  m_1182_io_x3; // @[MUL.scala 102:19]
  wire  m_1182_io_s; // @[MUL.scala 102:19]
  wire  m_1182_io_cout; // @[MUL.scala 102:19]
  wire  m_1183_io_x1; // @[MUL.scala 102:19]
  wire  m_1183_io_x2; // @[MUL.scala 102:19]
  wire  m_1183_io_x3; // @[MUL.scala 102:19]
  wire  m_1183_io_s; // @[MUL.scala 102:19]
  wire  m_1183_io_cout; // @[MUL.scala 102:19]
  wire  m_1184_io_x1; // @[MUL.scala 102:19]
  wire  m_1184_io_x2; // @[MUL.scala 102:19]
  wire  m_1184_io_x3; // @[MUL.scala 102:19]
  wire  m_1184_io_s; // @[MUL.scala 102:19]
  wire  m_1184_io_cout; // @[MUL.scala 102:19]
  wire  m_1185_io_x1; // @[MUL.scala 102:19]
  wire  m_1185_io_x2; // @[MUL.scala 102:19]
  wire  m_1185_io_x3; // @[MUL.scala 102:19]
  wire  m_1185_io_s; // @[MUL.scala 102:19]
  wire  m_1185_io_cout; // @[MUL.scala 102:19]
  wire  m_1186_io_x1; // @[MUL.scala 102:19]
  wire  m_1186_io_x2; // @[MUL.scala 102:19]
  wire  m_1186_io_x3; // @[MUL.scala 102:19]
  wire  m_1186_io_s; // @[MUL.scala 102:19]
  wire  m_1186_io_cout; // @[MUL.scala 102:19]
  wire  m_1187_io_in_0; // @[MUL.scala 124:19]
  wire  m_1187_io_in_1; // @[MUL.scala 124:19]
  wire  m_1187_io_out_0; // @[MUL.scala 124:19]
  wire  m_1187_io_out_1; // @[MUL.scala 124:19]
  wire  m_1188_io_x1; // @[MUL.scala 102:19]
  wire  m_1188_io_x2; // @[MUL.scala 102:19]
  wire  m_1188_io_x3; // @[MUL.scala 102:19]
  wire  m_1188_io_s; // @[MUL.scala 102:19]
  wire  m_1188_io_cout; // @[MUL.scala 102:19]
  wire  m_1189_io_x1; // @[MUL.scala 102:19]
  wire  m_1189_io_x2; // @[MUL.scala 102:19]
  wire  m_1189_io_x3; // @[MUL.scala 102:19]
  wire  m_1189_io_s; // @[MUL.scala 102:19]
  wire  m_1189_io_cout; // @[MUL.scala 102:19]
  wire  m_1190_io_x1; // @[MUL.scala 102:19]
  wire  m_1190_io_x2; // @[MUL.scala 102:19]
  wire  m_1190_io_x3; // @[MUL.scala 102:19]
  wire  m_1190_io_s; // @[MUL.scala 102:19]
  wire  m_1190_io_cout; // @[MUL.scala 102:19]
  wire  m_1191_io_x1; // @[MUL.scala 102:19]
  wire  m_1191_io_x2; // @[MUL.scala 102:19]
  wire  m_1191_io_x3; // @[MUL.scala 102:19]
  wire  m_1191_io_s; // @[MUL.scala 102:19]
  wire  m_1191_io_cout; // @[MUL.scala 102:19]
  wire  m_1192_io_x1; // @[MUL.scala 102:19]
  wire  m_1192_io_x2; // @[MUL.scala 102:19]
  wire  m_1192_io_x3; // @[MUL.scala 102:19]
  wire  m_1192_io_s; // @[MUL.scala 102:19]
  wire  m_1192_io_cout; // @[MUL.scala 102:19]
  wire  m_1193_io_x1; // @[MUL.scala 102:19]
  wire  m_1193_io_x2; // @[MUL.scala 102:19]
  wire  m_1193_io_x3; // @[MUL.scala 102:19]
  wire  m_1193_io_s; // @[MUL.scala 102:19]
  wire  m_1193_io_cout; // @[MUL.scala 102:19]
  wire  m_1194_io_x1; // @[MUL.scala 102:19]
  wire  m_1194_io_x2; // @[MUL.scala 102:19]
  wire  m_1194_io_x3; // @[MUL.scala 102:19]
  wire  m_1194_io_s; // @[MUL.scala 102:19]
  wire  m_1194_io_cout; // @[MUL.scala 102:19]
  wire  m_1195_io_x1; // @[MUL.scala 102:19]
  wire  m_1195_io_x2; // @[MUL.scala 102:19]
  wire  m_1195_io_x3; // @[MUL.scala 102:19]
  wire  m_1195_io_s; // @[MUL.scala 102:19]
  wire  m_1195_io_cout; // @[MUL.scala 102:19]
  wire  m_1196_io_x1; // @[MUL.scala 102:19]
  wire  m_1196_io_x2; // @[MUL.scala 102:19]
  wire  m_1196_io_x3; // @[MUL.scala 102:19]
  wire  m_1196_io_s; // @[MUL.scala 102:19]
  wire  m_1196_io_cout; // @[MUL.scala 102:19]
  wire  m_1197_io_x1; // @[MUL.scala 102:19]
  wire  m_1197_io_x2; // @[MUL.scala 102:19]
  wire  m_1197_io_x3; // @[MUL.scala 102:19]
  wire  m_1197_io_s; // @[MUL.scala 102:19]
  wire  m_1197_io_cout; // @[MUL.scala 102:19]
  wire  m_1198_io_x1; // @[MUL.scala 102:19]
  wire  m_1198_io_x2; // @[MUL.scala 102:19]
  wire  m_1198_io_x3; // @[MUL.scala 102:19]
  wire  m_1198_io_s; // @[MUL.scala 102:19]
  wire  m_1198_io_cout; // @[MUL.scala 102:19]
  wire  m_1199_io_x1; // @[MUL.scala 102:19]
  wire  m_1199_io_x2; // @[MUL.scala 102:19]
  wire  m_1199_io_x3; // @[MUL.scala 102:19]
  wire  m_1199_io_s; // @[MUL.scala 102:19]
  wire  m_1199_io_cout; // @[MUL.scala 102:19]
  wire  m_1200_io_x1; // @[MUL.scala 102:19]
  wire  m_1200_io_x2; // @[MUL.scala 102:19]
  wire  m_1200_io_x3; // @[MUL.scala 102:19]
  wire  m_1200_io_s; // @[MUL.scala 102:19]
  wire  m_1200_io_cout; // @[MUL.scala 102:19]
  wire  m_1201_io_x1; // @[MUL.scala 102:19]
  wire  m_1201_io_x2; // @[MUL.scala 102:19]
  wire  m_1201_io_x3; // @[MUL.scala 102:19]
  wire  m_1201_io_s; // @[MUL.scala 102:19]
  wire  m_1201_io_cout; // @[MUL.scala 102:19]
  wire  m_1202_io_x1; // @[MUL.scala 102:19]
  wire  m_1202_io_x2; // @[MUL.scala 102:19]
  wire  m_1202_io_x3; // @[MUL.scala 102:19]
  wire  m_1202_io_s; // @[MUL.scala 102:19]
  wire  m_1202_io_cout; // @[MUL.scala 102:19]
  wire  m_1203_io_x1; // @[MUL.scala 102:19]
  wire  m_1203_io_x2; // @[MUL.scala 102:19]
  wire  m_1203_io_x3; // @[MUL.scala 102:19]
  wire  m_1203_io_s; // @[MUL.scala 102:19]
  wire  m_1203_io_cout; // @[MUL.scala 102:19]
  wire  m_1204_io_x1; // @[MUL.scala 102:19]
  wire  m_1204_io_x2; // @[MUL.scala 102:19]
  wire  m_1204_io_x3; // @[MUL.scala 102:19]
  wire  m_1204_io_s; // @[MUL.scala 102:19]
  wire  m_1204_io_cout; // @[MUL.scala 102:19]
  wire  m_1205_io_x1; // @[MUL.scala 102:19]
  wire  m_1205_io_x2; // @[MUL.scala 102:19]
  wire  m_1205_io_x3; // @[MUL.scala 102:19]
  wire  m_1205_io_s; // @[MUL.scala 102:19]
  wire  m_1205_io_cout; // @[MUL.scala 102:19]
  wire  m_1206_io_x1; // @[MUL.scala 102:19]
  wire  m_1206_io_x2; // @[MUL.scala 102:19]
  wire  m_1206_io_x3; // @[MUL.scala 102:19]
  wire  m_1206_io_s; // @[MUL.scala 102:19]
  wire  m_1206_io_cout; // @[MUL.scala 102:19]
  wire  m_1207_io_x1; // @[MUL.scala 102:19]
  wire  m_1207_io_x2; // @[MUL.scala 102:19]
  wire  m_1207_io_x3; // @[MUL.scala 102:19]
  wire  m_1207_io_s; // @[MUL.scala 102:19]
  wire  m_1207_io_cout; // @[MUL.scala 102:19]
  wire  m_1208_io_x1; // @[MUL.scala 102:19]
  wire  m_1208_io_x2; // @[MUL.scala 102:19]
  wire  m_1208_io_x3; // @[MUL.scala 102:19]
  wire  m_1208_io_s; // @[MUL.scala 102:19]
  wire  m_1208_io_cout; // @[MUL.scala 102:19]
  wire  m_1209_io_x1; // @[MUL.scala 102:19]
  wire  m_1209_io_x2; // @[MUL.scala 102:19]
  wire  m_1209_io_x3; // @[MUL.scala 102:19]
  wire  m_1209_io_s; // @[MUL.scala 102:19]
  wire  m_1209_io_cout; // @[MUL.scala 102:19]
  wire  m_1210_io_x1; // @[MUL.scala 102:19]
  wire  m_1210_io_x2; // @[MUL.scala 102:19]
  wire  m_1210_io_x3; // @[MUL.scala 102:19]
  wire  m_1210_io_s; // @[MUL.scala 102:19]
  wire  m_1210_io_cout; // @[MUL.scala 102:19]
  wire  m_1211_io_x1; // @[MUL.scala 102:19]
  wire  m_1211_io_x2; // @[MUL.scala 102:19]
  wire  m_1211_io_x3; // @[MUL.scala 102:19]
  wire  m_1211_io_s; // @[MUL.scala 102:19]
  wire  m_1211_io_cout; // @[MUL.scala 102:19]
  wire  m_1212_io_x1; // @[MUL.scala 102:19]
  wire  m_1212_io_x2; // @[MUL.scala 102:19]
  wire  m_1212_io_x3; // @[MUL.scala 102:19]
  wire  m_1212_io_s; // @[MUL.scala 102:19]
  wire  m_1212_io_cout; // @[MUL.scala 102:19]
  wire  m_1213_io_x1; // @[MUL.scala 102:19]
  wire  m_1213_io_x2; // @[MUL.scala 102:19]
  wire  m_1213_io_x3; // @[MUL.scala 102:19]
  wire  m_1213_io_s; // @[MUL.scala 102:19]
  wire  m_1213_io_cout; // @[MUL.scala 102:19]
  wire  m_1214_io_x1; // @[MUL.scala 102:19]
  wire  m_1214_io_x2; // @[MUL.scala 102:19]
  wire  m_1214_io_x3; // @[MUL.scala 102:19]
  wire  m_1214_io_s; // @[MUL.scala 102:19]
  wire  m_1214_io_cout; // @[MUL.scala 102:19]
  wire  m_1215_io_x1; // @[MUL.scala 102:19]
  wire  m_1215_io_x2; // @[MUL.scala 102:19]
  wire  m_1215_io_x3; // @[MUL.scala 102:19]
  wire  m_1215_io_s; // @[MUL.scala 102:19]
  wire  m_1215_io_cout; // @[MUL.scala 102:19]
  wire  m_1216_io_x1; // @[MUL.scala 102:19]
  wire  m_1216_io_x2; // @[MUL.scala 102:19]
  wire  m_1216_io_x3; // @[MUL.scala 102:19]
  wire  m_1216_io_s; // @[MUL.scala 102:19]
  wire  m_1216_io_cout; // @[MUL.scala 102:19]
  wire  m_1217_io_x1; // @[MUL.scala 102:19]
  wire  m_1217_io_x2; // @[MUL.scala 102:19]
  wire  m_1217_io_x3; // @[MUL.scala 102:19]
  wire  m_1217_io_s; // @[MUL.scala 102:19]
  wire  m_1217_io_cout; // @[MUL.scala 102:19]
  wire  m_1218_io_x1; // @[MUL.scala 102:19]
  wire  m_1218_io_x2; // @[MUL.scala 102:19]
  wire  m_1218_io_x3; // @[MUL.scala 102:19]
  wire  m_1218_io_s; // @[MUL.scala 102:19]
  wire  m_1218_io_cout; // @[MUL.scala 102:19]
  wire  m_1219_io_x1; // @[MUL.scala 102:19]
  wire  m_1219_io_x2; // @[MUL.scala 102:19]
  wire  m_1219_io_x3; // @[MUL.scala 102:19]
  wire  m_1219_io_s; // @[MUL.scala 102:19]
  wire  m_1219_io_cout; // @[MUL.scala 102:19]
  wire  m_1220_io_x1; // @[MUL.scala 102:19]
  wire  m_1220_io_x2; // @[MUL.scala 102:19]
  wire  m_1220_io_x3; // @[MUL.scala 102:19]
  wire  m_1220_io_s; // @[MUL.scala 102:19]
  wire  m_1220_io_cout; // @[MUL.scala 102:19]
  wire  m_1221_io_x1; // @[MUL.scala 102:19]
  wire  m_1221_io_x2; // @[MUL.scala 102:19]
  wire  m_1221_io_x3; // @[MUL.scala 102:19]
  wire  m_1221_io_s; // @[MUL.scala 102:19]
  wire  m_1221_io_cout; // @[MUL.scala 102:19]
  wire  m_1222_io_in_0; // @[MUL.scala 124:19]
  wire  m_1222_io_in_1; // @[MUL.scala 124:19]
  wire  m_1222_io_out_0; // @[MUL.scala 124:19]
  wire  m_1222_io_out_1; // @[MUL.scala 124:19]
  wire  m_1223_io_x1; // @[MUL.scala 102:19]
  wire  m_1223_io_x2; // @[MUL.scala 102:19]
  wire  m_1223_io_x3; // @[MUL.scala 102:19]
  wire  m_1223_io_s; // @[MUL.scala 102:19]
  wire  m_1223_io_cout; // @[MUL.scala 102:19]
  wire  m_1224_io_x1; // @[MUL.scala 102:19]
  wire  m_1224_io_x2; // @[MUL.scala 102:19]
  wire  m_1224_io_x3; // @[MUL.scala 102:19]
  wire  m_1224_io_s; // @[MUL.scala 102:19]
  wire  m_1224_io_cout; // @[MUL.scala 102:19]
  wire  m_1225_io_x1; // @[MUL.scala 102:19]
  wire  m_1225_io_x2; // @[MUL.scala 102:19]
  wire  m_1225_io_x3; // @[MUL.scala 102:19]
  wire  m_1225_io_s; // @[MUL.scala 102:19]
  wire  m_1225_io_cout; // @[MUL.scala 102:19]
  wire  m_1226_io_x1; // @[MUL.scala 102:19]
  wire  m_1226_io_x2; // @[MUL.scala 102:19]
  wire  m_1226_io_x3; // @[MUL.scala 102:19]
  wire  m_1226_io_s; // @[MUL.scala 102:19]
  wire  m_1226_io_cout; // @[MUL.scala 102:19]
  wire  m_1227_io_in_0; // @[MUL.scala 124:19]
  wire  m_1227_io_in_1; // @[MUL.scala 124:19]
  wire  m_1227_io_out_0; // @[MUL.scala 124:19]
  wire  m_1227_io_out_1; // @[MUL.scala 124:19]
  wire  m_1228_io_x1; // @[MUL.scala 102:19]
  wire  m_1228_io_x2; // @[MUL.scala 102:19]
  wire  m_1228_io_x3; // @[MUL.scala 102:19]
  wire  m_1228_io_s; // @[MUL.scala 102:19]
  wire  m_1228_io_cout; // @[MUL.scala 102:19]
  wire  m_1229_io_x1; // @[MUL.scala 102:19]
  wire  m_1229_io_x2; // @[MUL.scala 102:19]
  wire  m_1229_io_x3; // @[MUL.scala 102:19]
  wire  m_1229_io_s; // @[MUL.scala 102:19]
  wire  m_1229_io_cout; // @[MUL.scala 102:19]
  wire  m_1230_io_x1; // @[MUL.scala 102:19]
  wire  m_1230_io_x2; // @[MUL.scala 102:19]
  wire  m_1230_io_x3; // @[MUL.scala 102:19]
  wire  m_1230_io_s; // @[MUL.scala 102:19]
  wire  m_1230_io_cout; // @[MUL.scala 102:19]
  wire  m_1231_io_x1; // @[MUL.scala 102:19]
  wire  m_1231_io_x2; // @[MUL.scala 102:19]
  wire  m_1231_io_x3; // @[MUL.scala 102:19]
  wire  m_1231_io_s; // @[MUL.scala 102:19]
  wire  m_1231_io_cout; // @[MUL.scala 102:19]
  wire  m_1232_io_in_0; // @[MUL.scala 124:19]
  wire  m_1232_io_in_1; // @[MUL.scala 124:19]
  wire  m_1232_io_out_0; // @[MUL.scala 124:19]
  wire  m_1232_io_out_1; // @[MUL.scala 124:19]
  wire  m_1233_io_x1; // @[MUL.scala 102:19]
  wire  m_1233_io_x2; // @[MUL.scala 102:19]
  wire  m_1233_io_x3; // @[MUL.scala 102:19]
  wire  m_1233_io_s; // @[MUL.scala 102:19]
  wire  m_1233_io_cout; // @[MUL.scala 102:19]
  wire  m_1234_io_x1; // @[MUL.scala 102:19]
  wire  m_1234_io_x2; // @[MUL.scala 102:19]
  wire  m_1234_io_x3; // @[MUL.scala 102:19]
  wire  m_1234_io_s; // @[MUL.scala 102:19]
  wire  m_1234_io_cout; // @[MUL.scala 102:19]
  wire  m_1235_io_x1; // @[MUL.scala 102:19]
  wire  m_1235_io_x2; // @[MUL.scala 102:19]
  wire  m_1235_io_x3; // @[MUL.scala 102:19]
  wire  m_1235_io_s; // @[MUL.scala 102:19]
  wire  m_1235_io_cout; // @[MUL.scala 102:19]
  wire  m_1236_io_x1; // @[MUL.scala 102:19]
  wire  m_1236_io_x2; // @[MUL.scala 102:19]
  wire  m_1236_io_x3; // @[MUL.scala 102:19]
  wire  m_1236_io_s; // @[MUL.scala 102:19]
  wire  m_1236_io_cout; // @[MUL.scala 102:19]
  wire  m_1237_io_in_0; // @[MUL.scala 124:19]
  wire  m_1237_io_in_1; // @[MUL.scala 124:19]
  wire  m_1237_io_out_0; // @[MUL.scala 124:19]
  wire  m_1237_io_out_1; // @[MUL.scala 124:19]
  wire  m_1238_io_x1; // @[MUL.scala 102:19]
  wire  m_1238_io_x2; // @[MUL.scala 102:19]
  wire  m_1238_io_x3; // @[MUL.scala 102:19]
  wire  m_1238_io_s; // @[MUL.scala 102:19]
  wire  m_1238_io_cout; // @[MUL.scala 102:19]
  wire  m_1239_io_x1; // @[MUL.scala 102:19]
  wire  m_1239_io_x2; // @[MUL.scala 102:19]
  wire  m_1239_io_x3; // @[MUL.scala 102:19]
  wire  m_1239_io_s; // @[MUL.scala 102:19]
  wire  m_1239_io_cout; // @[MUL.scala 102:19]
  wire  m_1240_io_x1; // @[MUL.scala 102:19]
  wire  m_1240_io_x2; // @[MUL.scala 102:19]
  wire  m_1240_io_x3; // @[MUL.scala 102:19]
  wire  m_1240_io_s; // @[MUL.scala 102:19]
  wire  m_1240_io_cout; // @[MUL.scala 102:19]
  wire  m_1241_io_x1; // @[MUL.scala 102:19]
  wire  m_1241_io_x2; // @[MUL.scala 102:19]
  wire  m_1241_io_x3; // @[MUL.scala 102:19]
  wire  m_1241_io_s; // @[MUL.scala 102:19]
  wire  m_1241_io_cout; // @[MUL.scala 102:19]
  wire  m_1242_io_in_0; // @[MUL.scala 124:19]
  wire  m_1242_io_in_1; // @[MUL.scala 124:19]
  wire  m_1242_io_out_0; // @[MUL.scala 124:19]
  wire  m_1242_io_out_1; // @[MUL.scala 124:19]
  wire  m_1243_io_x1; // @[MUL.scala 102:19]
  wire  m_1243_io_x2; // @[MUL.scala 102:19]
  wire  m_1243_io_x3; // @[MUL.scala 102:19]
  wire  m_1243_io_s; // @[MUL.scala 102:19]
  wire  m_1243_io_cout; // @[MUL.scala 102:19]
  wire  m_1244_io_x1; // @[MUL.scala 102:19]
  wire  m_1244_io_x2; // @[MUL.scala 102:19]
  wire  m_1244_io_x3; // @[MUL.scala 102:19]
  wire  m_1244_io_s; // @[MUL.scala 102:19]
  wire  m_1244_io_cout; // @[MUL.scala 102:19]
  wire  m_1245_io_x1; // @[MUL.scala 102:19]
  wire  m_1245_io_x2; // @[MUL.scala 102:19]
  wire  m_1245_io_x3; // @[MUL.scala 102:19]
  wire  m_1245_io_s; // @[MUL.scala 102:19]
  wire  m_1245_io_cout; // @[MUL.scala 102:19]
  wire  m_1246_io_x1; // @[MUL.scala 102:19]
  wire  m_1246_io_x2; // @[MUL.scala 102:19]
  wire  m_1246_io_x3; // @[MUL.scala 102:19]
  wire  m_1246_io_s; // @[MUL.scala 102:19]
  wire  m_1246_io_cout; // @[MUL.scala 102:19]
  wire  m_1247_io_x1; // @[MUL.scala 102:19]
  wire  m_1247_io_x2; // @[MUL.scala 102:19]
  wire  m_1247_io_x3; // @[MUL.scala 102:19]
  wire  m_1247_io_s; // @[MUL.scala 102:19]
  wire  m_1247_io_cout; // @[MUL.scala 102:19]
  wire  m_1248_io_x1; // @[MUL.scala 102:19]
  wire  m_1248_io_x2; // @[MUL.scala 102:19]
  wire  m_1248_io_x3; // @[MUL.scala 102:19]
  wire  m_1248_io_s; // @[MUL.scala 102:19]
  wire  m_1248_io_cout; // @[MUL.scala 102:19]
  wire  m_1249_io_x1; // @[MUL.scala 102:19]
  wire  m_1249_io_x2; // @[MUL.scala 102:19]
  wire  m_1249_io_x3; // @[MUL.scala 102:19]
  wire  m_1249_io_s; // @[MUL.scala 102:19]
  wire  m_1249_io_cout; // @[MUL.scala 102:19]
  wire  m_1250_io_x1; // @[MUL.scala 102:19]
  wire  m_1250_io_x2; // @[MUL.scala 102:19]
  wire  m_1250_io_x3; // @[MUL.scala 102:19]
  wire  m_1250_io_s; // @[MUL.scala 102:19]
  wire  m_1250_io_cout; // @[MUL.scala 102:19]
  wire  m_1251_io_x1; // @[MUL.scala 102:19]
  wire  m_1251_io_x2; // @[MUL.scala 102:19]
  wire  m_1251_io_x3; // @[MUL.scala 102:19]
  wire  m_1251_io_s; // @[MUL.scala 102:19]
  wire  m_1251_io_cout; // @[MUL.scala 102:19]
  wire  m_1252_io_x1; // @[MUL.scala 102:19]
  wire  m_1252_io_x2; // @[MUL.scala 102:19]
  wire  m_1252_io_x3; // @[MUL.scala 102:19]
  wire  m_1252_io_s; // @[MUL.scala 102:19]
  wire  m_1252_io_cout; // @[MUL.scala 102:19]
  wire  m_1253_io_x1; // @[MUL.scala 102:19]
  wire  m_1253_io_x2; // @[MUL.scala 102:19]
  wire  m_1253_io_x3; // @[MUL.scala 102:19]
  wire  m_1253_io_s; // @[MUL.scala 102:19]
  wire  m_1253_io_cout; // @[MUL.scala 102:19]
  wire  m_1254_io_x1; // @[MUL.scala 102:19]
  wire  m_1254_io_x2; // @[MUL.scala 102:19]
  wire  m_1254_io_x3; // @[MUL.scala 102:19]
  wire  m_1254_io_s; // @[MUL.scala 102:19]
  wire  m_1254_io_cout; // @[MUL.scala 102:19]
  wire  m_1255_io_x1; // @[MUL.scala 102:19]
  wire  m_1255_io_x2; // @[MUL.scala 102:19]
  wire  m_1255_io_x3; // @[MUL.scala 102:19]
  wire  m_1255_io_s; // @[MUL.scala 102:19]
  wire  m_1255_io_cout; // @[MUL.scala 102:19]
  wire  m_1256_io_x1; // @[MUL.scala 102:19]
  wire  m_1256_io_x2; // @[MUL.scala 102:19]
  wire  m_1256_io_x3; // @[MUL.scala 102:19]
  wire  m_1256_io_s; // @[MUL.scala 102:19]
  wire  m_1256_io_cout; // @[MUL.scala 102:19]
  wire  m_1257_io_x1; // @[MUL.scala 102:19]
  wire  m_1257_io_x2; // @[MUL.scala 102:19]
  wire  m_1257_io_x3; // @[MUL.scala 102:19]
  wire  m_1257_io_s; // @[MUL.scala 102:19]
  wire  m_1257_io_cout; // @[MUL.scala 102:19]
  wire  m_1258_io_x1; // @[MUL.scala 102:19]
  wire  m_1258_io_x2; // @[MUL.scala 102:19]
  wire  m_1258_io_x3; // @[MUL.scala 102:19]
  wire  m_1258_io_s; // @[MUL.scala 102:19]
  wire  m_1258_io_cout; // @[MUL.scala 102:19]
  wire  m_1259_io_x1; // @[MUL.scala 102:19]
  wire  m_1259_io_x2; // @[MUL.scala 102:19]
  wire  m_1259_io_x3; // @[MUL.scala 102:19]
  wire  m_1259_io_s; // @[MUL.scala 102:19]
  wire  m_1259_io_cout; // @[MUL.scala 102:19]
  wire  m_1260_io_x1; // @[MUL.scala 102:19]
  wire  m_1260_io_x2; // @[MUL.scala 102:19]
  wire  m_1260_io_x3; // @[MUL.scala 102:19]
  wire  m_1260_io_s; // @[MUL.scala 102:19]
  wire  m_1260_io_cout; // @[MUL.scala 102:19]
  wire  m_1261_io_x1; // @[MUL.scala 102:19]
  wire  m_1261_io_x2; // @[MUL.scala 102:19]
  wire  m_1261_io_x3; // @[MUL.scala 102:19]
  wire  m_1261_io_s; // @[MUL.scala 102:19]
  wire  m_1261_io_cout; // @[MUL.scala 102:19]
  wire  m_1262_io_x1; // @[MUL.scala 102:19]
  wire  m_1262_io_x2; // @[MUL.scala 102:19]
  wire  m_1262_io_x3; // @[MUL.scala 102:19]
  wire  m_1262_io_s; // @[MUL.scala 102:19]
  wire  m_1262_io_cout; // @[MUL.scala 102:19]
  wire  m_1263_io_x1; // @[MUL.scala 102:19]
  wire  m_1263_io_x2; // @[MUL.scala 102:19]
  wire  m_1263_io_x3; // @[MUL.scala 102:19]
  wire  m_1263_io_s; // @[MUL.scala 102:19]
  wire  m_1263_io_cout; // @[MUL.scala 102:19]
  wire  m_1264_io_x1; // @[MUL.scala 102:19]
  wire  m_1264_io_x2; // @[MUL.scala 102:19]
  wire  m_1264_io_x3; // @[MUL.scala 102:19]
  wire  m_1264_io_s; // @[MUL.scala 102:19]
  wire  m_1264_io_cout; // @[MUL.scala 102:19]
  wire  m_1265_io_x1; // @[MUL.scala 102:19]
  wire  m_1265_io_x2; // @[MUL.scala 102:19]
  wire  m_1265_io_x3; // @[MUL.scala 102:19]
  wire  m_1265_io_s; // @[MUL.scala 102:19]
  wire  m_1265_io_cout; // @[MUL.scala 102:19]
  wire  m_1266_io_x1; // @[MUL.scala 102:19]
  wire  m_1266_io_x2; // @[MUL.scala 102:19]
  wire  m_1266_io_x3; // @[MUL.scala 102:19]
  wire  m_1266_io_s; // @[MUL.scala 102:19]
  wire  m_1266_io_cout; // @[MUL.scala 102:19]
  wire  m_1267_io_x1; // @[MUL.scala 102:19]
  wire  m_1267_io_x2; // @[MUL.scala 102:19]
  wire  m_1267_io_x3; // @[MUL.scala 102:19]
  wire  m_1267_io_s; // @[MUL.scala 102:19]
  wire  m_1267_io_cout; // @[MUL.scala 102:19]
  wire  m_1268_io_x1; // @[MUL.scala 102:19]
  wire  m_1268_io_x2; // @[MUL.scala 102:19]
  wire  m_1268_io_x3; // @[MUL.scala 102:19]
  wire  m_1268_io_s; // @[MUL.scala 102:19]
  wire  m_1268_io_cout; // @[MUL.scala 102:19]
  wire  m_1269_io_x1; // @[MUL.scala 102:19]
  wire  m_1269_io_x2; // @[MUL.scala 102:19]
  wire  m_1269_io_x3; // @[MUL.scala 102:19]
  wire  m_1269_io_s; // @[MUL.scala 102:19]
  wire  m_1269_io_cout; // @[MUL.scala 102:19]
  wire  m_1270_io_in_0; // @[MUL.scala 124:19]
  wire  m_1270_io_in_1; // @[MUL.scala 124:19]
  wire  m_1270_io_out_0; // @[MUL.scala 124:19]
  wire  m_1270_io_out_1; // @[MUL.scala 124:19]
  wire  m_1271_io_x1; // @[MUL.scala 102:19]
  wire  m_1271_io_x2; // @[MUL.scala 102:19]
  wire  m_1271_io_x3; // @[MUL.scala 102:19]
  wire  m_1271_io_s; // @[MUL.scala 102:19]
  wire  m_1271_io_cout; // @[MUL.scala 102:19]
  wire  m_1272_io_x1; // @[MUL.scala 102:19]
  wire  m_1272_io_x2; // @[MUL.scala 102:19]
  wire  m_1272_io_x3; // @[MUL.scala 102:19]
  wire  m_1272_io_s; // @[MUL.scala 102:19]
  wire  m_1272_io_cout; // @[MUL.scala 102:19]
  wire  m_1273_io_x1; // @[MUL.scala 102:19]
  wire  m_1273_io_x2; // @[MUL.scala 102:19]
  wire  m_1273_io_x3; // @[MUL.scala 102:19]
  wire  m_1273_io_s; // @[MUL.scala 102:19]
  wire  m_1273_io_cout; // @[MUL.scala 102:19]
  wire  m_1274_io_x1; // @[MUL.scala 102:19]
  wire  m_1274_io_x2; // @[MUL.scala 102:19]
  wire  m_1274_io_x3; // @[MUL.scala 102:19]
  wire  m_1274_io_s; // @[MUL.scala 102:19]
  wire  m_1274_io_cout; // @[MUL.scala 102:19]
  wire  m_1275_io_x1; // @[MUL.scala 102:19]
  wire  m_1275_io_x2; // @[MUL.scala 102:19]
  wire  m_1275_io_x3; // @[MUL.scala 102:19]
  wire  m_1275_io_s; // @[MUL.scala 102:19]
  wire  m_1275_io_cout; // @[MUL.scala 102:19]
  wire  m_1276_io_x1; // @[MUL.scala 102:19]
  wire  m_1276_io_x2; // @[MUL.scala 102:19]
  wire  m_1276_io_x3; // @[MUL.scala 102:19]
  wire  m_1276_io_s; // @[MUL.scala 102:19]
  wire  m_1276_io_cout; // @[MUL.scala 102:19]
  wire  m_1277_io_x1; // @[MUL.scala 102:19]
  wire  m_1277_io_x2; // @[MUL.scala 102:19]
  wire  m_1277_io_x3; // @[MUL.scala 102:19]
  wire  m_1277_io_s; // @[MUL.scala 102:19]
  wire  m_1277_io_cout; // @[MUL.scala 102:19]
  wire  m_1278_io_x1; // @[MUL.scala 102:19]
  wire  m_1278_io_x2; // @[MUL.scala 102:19]
  wire  m_1278_io_x3; // @[MUL.scala 102:19]
  wire  m_1278_io_s; // @[MUL.scala 102:19]
  wire  m_1278_io_cout; // @[MUL.scala 102:19]
  wire  m_1279_io_x1; // @[MUL.scala 102:19]
  wire  m_1279_io_x2; // @[MUL.scala 102:19]
  wire  m_1279_io_x3; // @[MUL.scala 102:19]
  wire  m_1279_io_s; // @[MUL.scala 102:19]
  wire  m_1279_io_cout; // @[MUL.scala 102:19]
  wire  m_1280_io_x1; // @[MUL.scala 102:19]
  wire  m_1280_io_x2; // @[MUL.scala 102:19]
  wire  m_1280_io_x3; // @[MUL.scala 102:19]
  wire  m_1280_io_s; // @[MUL.scala 102:19]
  wire  m_1280_io_cout; // @[MUL.scala 102:19]
  wire  m_1281_io_x1; // @[MUL.scala 102:19]
  wire  m_1281_io_x2; // @[MUL.scala 102:19]
  wire  m_1281_io_x3; // @[MUL.scala 102:19]
  wire  m_1281_io_s; // @[MUL.scala 102:19]
  wire  m_1281_io_cout; // @[MUL.scala 102:19]
  wire  m_1282_io_x1; // @[MUL.scala 102:19]
  wire  m_1282_io_x2; // @[MUL.scala 102:19]
  wire  m_1282_io_x3; // @[MUL.scala 102:19]
  wire  m_1282_io_s; // @[MUL.scala 102:19]
  wire  m_1282_io_cout; // @[MUL.scala 102:19]
  wire  m_1283_io_x1; // @[MUL.scala 102:19]
  wire  m_1283_io_x2; // @[MUL.scala 102:19]
  wire  m_1283_io_x3; // @[MUL.scala 102:19]
  wire  m_1283_io_s; // @[MUL.scala 102:19]
  wire  m_1283_io_cout; // @[MUL.scala 102:19]
  wire  m_1284_io_x1; // @[MUL.scala 102:19]
  wire  m_1284_io_x2; // @[MUL.scala 102:19]
  wire  m_1284_io_x3; // @[MUL.scala 102:19]
  wire  m_1284_io_s; // @[MUL.scala 102:19]
  wire  m_1284_io_cout; // @[MUL.scala 102:19]
  wire  m_1285_io_x1; // @[MUL.scala 102:19]
  wire  m_1285_io_x2; // @[MUL.scala 102:19]
  wire  m_1285_io_x3; // @[MUL.scala 102:19]
  wire  m_1285_io_s; // @[MUL.scala 102:19]
  wire  m_1285_io_cout; // @[MUL.scala 102:19]
  wire  m_1286_io_x1; // @[MUL.scala 102:19]
  wire  m_1286_io_x2; // @[MUL.scala 102:19]
  wire  m_1286_io_x3; // @[MUL.scala 102:19]
  wire  m_1286_io_s; // @[MUL.scala 102:19]
  wire  m_1286_io_cout; // @[MUL.scala 102:19]
  wire  m_1287_io_x1; // @[MUL.scala 102:19]
  wire  m_1287_io_x2; // @[MUL.scala 102:19]
  wire  m_1287_io_x3; // @[MUL.scala 102:19]
  wire  m_1287_io_s; // @[MUL.scala 102:19]
  wire  m_1287_io_cout; // @[MUL.scala 102:19]
  wire  m_1288_io_x1; // @[MUL.scala 102:19]
  wire  m_1288_io_x2; // @[MUL.scala 102:19]
  wire  m_1288_io_x3; // @[MUL.scala 102:19]
  wire  m_1288_io_s; // @[MUL.scala 102:19]
  wire  m_1288_io_cout; // @[MUL.scala 102:19]
  wire  m_1289_io_x1; // @[MUL.scala 102:19]
  wire  m_1289_io_x2; // @[MUL.scala 102:19]
  wire  m_1289_io_x3; // @[MUL.scala 102:19]
  wire  m_1289_io_s; // @[MUL.scala 102:19]
  wire  m_1289_io_cout; // @[MUL.scala 102:19]
  wire  m_1290_io_x1; // @[MUL.scala 102:19]
  wire  m_1290_io_x2; // @[MUL.scala 102:19]
  wire  m_1290_io_x3; // @[MUL.scala 102:19]
  wire  m_1290_io_s; // @[MUL.scala 102:19]
  wire  m_1290_io_cout; // @[MUL.scala 102:19]
  wire  m_1291_io_in_0; // @[MUL.scala 124:19]
  wire  m_1291_io_in_1; // @[MUL.scala 124:19]
  wire  m_1291_io_out_0; // @[MUL.scala 124:19]
  wire  m_1291_io_out_1; // @[MUL.scala 124:19]
  wire  m_1292_io_x1; // @[MUL.scala 102:19]
  wire  m_1292_io_x2; // @[MUL.scala 102:19]
  wire  m_1292_io_x3; // @[MUL.scala 102:19]
  wire  m_1292_io_s; // @[MUL.scala 102:19]
  wire  m_1292_io_cout; // @[MUL.scala 102:19]
  wire  m_1293_io_x1; // @[MUL.scala 102:19]
  wire  m_1293_io_x2; // @[MUL.scala 102:19]
  wire  m_1293_io_x3; // @[MUL.scala 102:19]
  wire  m_1293_io_s; // @[MUL.scala 102:19]
  wire  m_1293_io_cout; // @[MUL.scala 102:19]
  wire  m_1294_io_in_0; // @[MUL.scala 124:19]
  wire  m_1294_io_in_1; // @[MUL.scala 124:19]
  wire  m_1294_io_out_0; // @[MUL.scala 124:19]
  wire  m_1294_io_out_1; // @[MUL.scala 124:19]
  wire  m_1295_io_x1; // @[MUL.scala 102:19]
  wire  m_1295_io_x2; // @[MUL.scala 102:19]
  wire  m_1295_io_x3; // @[MUL.scala 102:19]
  wire  m_1295_io_s; // @[MUL.scala 102:19]
  wire  m_1295_io_cout; // @[MUL.scala 102:19]
  wire  m_1296_io_x1; // @[MUL.scala 102:19]
  wire  m_1296_io_x2; // @[MUL.scala 102:19]
  wire  m_1296_io_x3; // @[MUL.scala 102:19]
  wire  m_1296_io_s; // @[MUL.scala 102:19]
  wire  m_1296_io_cout; // @[MUL.scala 102:19]
  wire  m_1297_io_in_0; // @[MUL.scala 124:19]
  wire  m_1297_io_in_1; // @[MUL.scala 124:19]
  wire  m_1297_io_out_0; // @[MUL.scala 124:19]
  wire  m_1297_io_out_1; // @[MUL.scala 124:19]
  wire  m_1298_io_x1; // @[MUL.scala 102:19]
  wire  m_1298_io_x2; // @[MUL.scala 102:19]
  wire  m_1298_io_x3; // @[MUL.scala 102:19]
  wire  m_1298_io_s; // @[MUL.scala 102:19]
  wire  m_1298_io_cout; // @[MUL.scala 102:19]
  wire  m_1299_io_x1; // @[MUL.scala 102:19]
  wire  m_1299_io_x2; // @[MUL.scala 102:19]
  wire  m_1299_io_x3; // @[MUL.scala 102:19]
  wire  m_1299_io_s; // @[MUL.scala 102:19]
  wire  m_1299_io_cout; // @[MUL.scala 102:19]
  wire  m_1300_io_in_0; // @[MUL.scala 124:19]
  wire  m_1300_io_in_1; // @[MUL.scala 124:19]
  wire  m_1300_io_out_0; // @[MUL.scala 124:19]
  wire  m_1300_io_out_1; // @[MUL.scala 124:19]
  wire  m_1301_io_x1; // @[MUL.scala 102:19]
  wire  m_1301_io_x2; // @[MUL.scala 102:19]
  wire  m_1301_io_x3; // @[MUL.scala 102:19]
  wire  m_1301_io_s; // @[MUL.scala 102:19]
  wire  m_1301_io_cout; // @[MUL.scala 102:19]
  wire  m_1302_io_x1; // @[MUL.scala 102:19]
  wire  m_1302_io_x2; // @[MUL.scala 102:19]
  wire  m_1302_io_x3; // @[MUL.scala 102:19]
  wire  m_1302_io_s; // @[MUL.scala 102:19]
  wire  m_1302_io_cout; // @[MUL.scala 102:19]
  wire  m_1303_io_in_0; // @[MUL.scala 124:19]
  wire  m_1303_io_in_1; // @[MUL.scala 124:19]
  wire  m_1303_io_out_0; // @[MUL.scala 124:19]
  wire  m_1303_io_out_1; // @[MUL.scala 124:19]
  wire  m_1304_io_x1; // @[MUL.scala 102:19]
  wire  m_1304_io_x2; // @[MUL.scala 102:19]
  wire  m_1304_io_x3; // @[MUL.scala 102:19]
  wire  m_1304_io_s; // @[MUL.scala 102:19]
  wire  m_1304_io_cout; // @[MUL.scala 102:19]
  wire  m_1305_io_x1; // @[MUL.scala 102:19]
  wire  m_1305_io_x2; // @[MUL.scala 102:19]
  wire  m_1305_io_x3; // @[MUL.scala 102:19]
  wire  m_1305_io_s; // @[MUL.scala 102:19]
  wire  m_1305_io_cout; // @[MUL.scala 102:19]
  wire  m_1306_io_x1; // @[MUL.scala 102:19]
  wire  m_1306_io_x2; // @[MUL.scala 102:19]
  wire  m_1306_io_x3; // @[MUL.scala 102:19]
  wire  m_1306_io_s; // @[MUL.scala 102:19]
  wire  m_1306_io_cout; // @[MUL.scala 102:19]
  wire  m_1307_io_x1; // @[MUL.scala 102:19]
  wire  m_1307_io_x2; // @[MUL.scala 102:19]
  wire  m_1307_io_x3; // @[MUL.scala 102:19]
  wire  m_1307_io_s; // @[MUL.scala 102:19]
  wire  m_1307_io_cout; // @[MUL.scala 102:19]
  wire  m_1308_io_x1; // @[MUL.scala 102:19]
  wire  m_1308_io_x2; // @[MUL.scala 102:19]
  wire  m_1308_io_x3; // @[MUL.scala 102:19]
  wire  m_1308_io_s; // @[MUL.scala 102:19]
  wire  m_1308_io_cout; // @[MUL.scala 102:19]
  wire  m_1309_io_x1; // @[MUL.scala 102:19]
  wire  m_1309_io_x2; // @[MUL.scala 102:19]
  wire  m_1309_io_x3; // @[MUL.scala 102:19]
  wire  m_1309_io_s; // @[MUL.scala 102:19]
  wire  m_1309_io_cout; // @[MUL.scala 102:19]
  wire  m_1310_io_x1; // @[MUL.scala 102:19]
  wire  m_1310_io_x2; // @[MUL.scala 102:19]
  wire  m_1310_io_x3; // @[MUL.scala 102:19]
  wire  m_1310_io_s; // @[MUL.scala 102:19]
  wire  m_1310_io_cout; // @[MUL.scala 102:19]
  wire  m_1311_io_x1; // @[MUL.scala 102:19]
  wire  m_1311_io_x2; // @[MUL.scala 102:19]
  wire  m_1311_io_x3; // @[MUL.scala 102:19]
  wire  m_1311_io_s; // @[MUL.scala 102:19]
  wire  m_1311_io_cout; // @[MUL.scala 102:19]
  wire  m_1312_io_x1; // @[MUL.scala 102:19]
  wire  m_1312_io_x2; // @[MUL.scala 102:19]
  wire  m_1312_io_x3; // @[MUL.scala 102:19]
  wire  m_1312_io_s; // @[MUL.scala 102:19]
  wire  m_1312_io_cout; // @[MUL.scala 102:19]
  wire  m_1313_io_x1; // @[MUL.scala 102:19]
  wire  m_1313_io_x2; // @[MUL.scala 102:19]
  wire  m_1313_io_x3; // @[MUL.scala 102:19]
  wire  m_1313_io_s; // @[MUL.scala 102:19]
  wire  m_1313_io_cout; // @[MUL.scala 102:19]
  wire  m_1314_io_x1; // @[MUL.scala 102:19]
  wire  m_1314_io_x2; // @[MUL.scala 102:19]
  wire  m_1314_io_x3; // @[MUL.scala 102:19]
  wire  m_1314_io_s; // @[MUL.scala 102:19]
  wire  m_1314_io_cout; // @[MUL.scala 102:19]
  wire  m_1315_io_x1; // @[MUL.scala 102:19]
  wire  m_1315_io_x2; // @[MUL.scala 102:19]
  wire  m_1315_io_x3; // @[MUL.scala 102:19]
  wire  m_1315_io_s; // @[MUL.scala 102:19]
  wire  m_1315_io_cout; // @[MUL.scala 102:19]
  wire  m_1316_io_x1; // @[MUL.scala 102:19]
  wire  m_1316_io_x2; // @[MUL.scala 102:19]
  wire  m_1316_io_x3; // @[MUL.scala 102:19]
  wire  m_1316_io_s; // @[MUL.scala 102:19]
  wire  m_1316_io_cout; // @[MUL.scala 102:19]
  wire  m_1317_io_in_0; // @[MUL.scala 124:19]
  wire  m_1317_io_in_1; // @[MUL.scala 124:19]
  wire  m_1317_io_out_0; // @[MUL.scala 124:19]
  wire  m_1317_io_out_1; // @[MUL.scala 124:19]
  wire  m_1318_io_x1; // @[MUL.scala 102:19]
  wire  m_1318_io_x2; // @[MUL.scala 102:19]
  wire  m_1318_io_x3; // @[MUL.scala 102:19]
  wire  m_1318_io_s; // @[MUL.scala 102:19]
  wire  m_1318_io_cout; // @[MUL.scala 102:19]
  wire  m_1319_io_x1; // @[MUL.scala 102:19]
  wire  m_1319_io_x2; // @[MUL.scala 102:19]
  wire  m_1319_io_x3; // @[MUL.scala 102:19]
  wire  m_1319_io_s; // @[MUL.scala 102:19]
  wire  m_1319_io_cout; // @[MUL.scala 102:19]
  wire  m_1320_io_x1; // @[MUL.scala 102:19]
  wire  m_1320_io_x2; // @[MUL.scala 102:19]
  wire  m_1320_io_x3; // @[MUL.scala 102:19]
  wire  m_1320_io_s; // @[MUL.scala 102:19]
  wire  m_1320_io_cout; // @[MUL.scala 102:19]
  wire  m_1321_io_x1; // @[MUL.scala 102:19]
  wire  m_1321_io_x2; // @[MUL.scala 102:19]
  wire  m_1321_io_x3; // @[MUL.scala 102:19]
  wire  m_1321_io_s; // @[MUL.scala 102:19]
  wire  m_1321_io_cout; // @[MUL.scala 102:19]
  wire  m_1322_io_x1; // @[MUL.scala 102:19]
  wire  m_1322_io_x2; // @[MUL.scala 102:19]
  wire  m_1322_io_x3; // @[MUL.scala 102:19]
  wire  m_1322_io_s; // @[MUL.scala 102:19]
  wire  m_1322_io_cout; // @[MUL.scala 102:19]
  wire  m_1323_io_x1; // @[MUL.scala 102:19]
  wire  m_1323_io_x2; // @[MUL.scala 102:19]
  wire  m_1323_io_x3; // @[MUL.scala 102:19]
  wire  m_1323_io_s; // @[MUL.scala 102:19]
  wire  m_1323_io_cout; // @[MUL.scala 102:19]
  wire  m_1324_io_in_0; // @[MUL.scala 124:19]
  wire  m_1324_io_in_1; // @[MUL.scala 124:19]
  wire  m_1324_io_out_0; // @[MUL.scala 124:19]
  wire  m_1324_io_out_1; // @[MUL.scala 124:19]
  wire  m_1325_io_in_0; // @[MUL.scala 124:19]
  wire  m_1325_io_in_1; // @[MUL.scala 124:19]
  wire  m_1325_io_out_0; // @[MUL.scala 124:19]
  wire  m_1325_io_out_1; // @[MUL.scala 124:19]
  wire  m_1326_io_in_0; // @[MUL.scala 124:19]
  wire  m_1326_io_in_1; // @[MUL.scala 124:19]
  wire  m_1326_io_out_0; // @[MUL.scala 124:19]
  wire  m_1326_io_out_1; // @[MUL.scala 124:19]
  wire  m_1327_io_in_0; // @[MUL.scala 124:19]
  wire  m_1327_io_in_1; // @[MUL.scala 124:19]
  wire  m_1327_io_out_0; // @[MUL.scala 124:19]
  wire  m_1327_io_out_1; // @[MUL.scala 124:19]
  wire  m_1328_io_in_0; // @[MUL.scala 124:19]
  wire  m_1328_io_in_1; // @[MUL.scala 124:19]
  wire  m_1328_io_out_0; // @[MUL.scala 124:19]
  wire  m_1328_io_out_1; // @[MUL.scala 124:19]
  wire  m_1329_io_in_0; // @[MUL.scala 124:19]
  wire  m_1329_io_in_1; // @[MUL.scala 124:19]
  wire  m_1329_io_out_0; // @[MUL.scala 124:19]
  wire  m_1329_io_out_1; // @[MUL.scala 124:19]
  wire  m_1330_io_in_0; // @[MUL.scala 124:19]
  wire  m_1330_io_in_1; // @[MUL.scala 124:19]
  wire  m_1330_io_out_0; // @[MUL.scala 124:19]
  wire  m_1330_io_out_1; // @[MUL.scala 124:19]
  wire  m_1331_io_in_0; // @[MUL.scala 124:19]
  wire  m_1331_io_in_1; // @[MUL.scala 124:19]
  wire  m_1331_io_out_0; // @[MUL.scala 124:19]
  wire  m_1331_io_out_1; // @[MUL.scala 124:19]
  wire  m_1332_io_in_0; // @[MUL.scala 124:19]
  wire  m_1332_io_in_1; // @[MUL.scala 124:19]
  wire  m_1332_io_out_0; // @[MUL.scala 124:19]
  wire  m_1332_io_out_1; // @[MUL.scala 124:19]
  wire  m_1333_io_in_0; // @[MUL.scala 124:19]
  wire  m_1333_io_in_1; // @[MUL.scala 124:19]
  wire  m_1333_io_out_0; // @[MUL.scala 124:19]
  wire  m_1333_io_out_1; // @[MUL.scala 124:19]
  wire  m_1334_io_x1; // @[MUL.scala 102:19]
  wire  m_1334_io_x2; // @[MUL.scala 102:19]
  wire  m_1334_io_x3; // @[MUL.scala 102:19]
  wire  m_1334_io_s; // @[MUL.scala 102:19]
  wire  m_1334_io_cout; // @[MUL.scala 102:19]
  wire  m_1335_io_x1; // @[MUL.scala 102:19]
  wire  m_1335_io_x2; // @[MUL.scala 102:19]
  wire  m_1335_io_x3; // @[MUL.scala 102:19]
  wire  m_1335_io_s; // @[MUL.scala 102:19]
  wire  m_1335_io_cout; // @[MUL.scala 102:19]
  wire  m_1336_io_x1; // @[MUL.scala 102:19]
  wire  m_1336_io_x2; // @[MUL.scala 102:19]
  wire  m_1336_io_x3; // @[MUL.scala 102:19]
  wire  m_1336_io_s; // @[MUL.scala 102:19]
  wire  m_1336_io_cout; // @[MUL.scala 102:19]
  wire  m_1337_io_x1; // @[MUL.scala 102:19]
  wire  m_1337_io_x2; // @[MUL.scala 102:19]
  wire  m_1337_io_x3; // @[MUL.scala 102:19]
  wire  m_1337_io_s; // @[MUL.scala 102:19]
  wire  m_1337_io_cout; // @[MUL.scala 102:19]
  wire  m_1338_io_x1; // @[MUL.scala 102:19]
  wire  m_1338_io_x2; // @[MUL.scala 102:19]
  wire  m_1338_io_x3; // @[MUL.scala 102:19]
  wire  m_1338_io_s; // @[MUL.scala 102:19]
  wire  m_1338_io_cout; // @[MUL.scala 102:19]
  wire  m_1339_io_x1; // @[MUL.scala 102:19]
  wire  m_1339_io_x2; // @[MUL.scala 102:19]
  wire  m_1339_io_x3; // @[MUL.scala 102:19]
  wire  m_1339_io_s; // @[MUL.scala 102:19]
  wire  m_1339_io_cout; // @[MUL.scala 102:19]
  wire  m_1340_io_x1; // @[MUL.scala 102:19]
  wire  m_1340_io_x2; // @[MUL.scala 102:19]
  wire  m_1340_io_x3; // @[MUL.scala 102:19]
  wire  m_1340_io_s; // @[MUL.scala 102:19]
  wire  m_1340_io_cout; // @[MUL.scala 102:19]
  wire  m_1341_io_x1; // @[MUL.scala 102:19]
  wire  m_1341_io_x2; // @[MUL.scala 102:19]
  wire  m_1341_io_x3; // @[MUL.scala 102:19]
  wire  m_1341_io_s; // @[MUL.scala 102:19]
  wire  m_1341_io_cout; // @[MUL.scala 102:19]
  wire  m_1342_io_x1; // @[MUL.scala 102:19]
  wire  m_1342_io_x2; // @[MUL.scala 102:19]
  wire  m_1342_io_x3; // @[MUL.scala 102:19]
  wire  m_1342_io_s; // @[MUL.scala 102:19]
  wire  m_1342_io_cout; // @[MUL.scala 102:19]
  wire  m_1343_io_x1; // @[MUL.scala 102:19]
  wire  m_1343_io_x2; // @[MUL.scala 102:19]
  wire  m_1343_io_x3; // @[MUL.scala 102:19]
  wire  m_1343_io_s; // @[MUL.scala 102:19]
  wire  m_1343_io_cout; // @[MUL.scala 102:19]
  wire  m_1344_io_in_0; // @[MUL.scala 124:19]
  wire  m_1344_io_in_1; // @[MUL.scala 124:19]
  wire  m_1344_io_out_0; // @[MUL.scala 124:19]
  wire  m_1344_io_out_1; // @[MUL.scala 124:19]
  wire  m_1345_io_x1; // @[MUL.scala 102:19]
  wire  m_1345_io_x2; // @[MUL.scala 102:19]
  wire  m_1345_io_x3; // @[MUL.scala 102:19]
  wire  m_1345_io_s; // @[MUL.scala 102:19]
  wire  m_1345_io_cout; // @[MUL.scala 102:19]
  wire  m_1346_io_in_0; // @[MUL.scala 124:19]
  wire  m_1346_io_in_1; // @[MUL.scala 124:19]
  wire  m_1346_io_out_0; // @[MUL.scala 124:19]
  wire  m_1346_io_out_1; // @[MUL.scala 124:19]
  wire  m_1347_io_x1; // @[MUL.scala 102:19]
  wire  m_1347_io_x2; // @[MUL.scala 102:19]
  wire  m_1347_io_x3; // @[MUL.scala 102:19]
  wire  m_1347_io_s; // @[MUL.scala 102:19]
  wire  m_1347_io_cout; // @[MUL.scala 102:19]
  wire  m_1348_io_in_0; // @[MUL.scala 124:19]
  wire  m_1348_io_in_1; // @[MUL.scala 124:19]
  wire  m_1348_io_out_0; // @[MUL.scala 124:19]
  wire  m_1348_io_out_1; // @[MUL.scala 124:19]
  wire  m_1349_io_x1; // @[MUL.scala 102:19]
  wire  m_1349_io_x2; // @[MUL.scala 102:19]
  wire  m_1349_io_x3; // @[MUL.scala 102:19]
  wire  m_1349_io_s; // @[MUL.scala 102:19]
  wire  m_1349_io_cout; // @[MUL.scala 102:19]
  wire  m_1350_io_in_0; // @[MUL.scala 124:19]
  wire  m_1350_io_in_1; // @[MUL.scala 124:19]
  wire  m_1350_io_out_0; // @[MUL.scala 124:19]
  wire  m_1350_io_out_1; // @[MUL.scala 124:19]
  wire  m_1351_io_x1; // @[MUL.scala 102:19]
  wire  m_1351_io_x2; // @[MUL.scala 102:19]
  wire  m_1351_io_x3; // @[MUL.scala 102:19]
  wire  m_1351_io_s; // @[MUL.scala 102:19]
  wire  m_1351_io_cout; // @[MUL.scala 102:19]
  wire  m_1352_io_x1; // @[MUL.scala 102:19]
  wire  m_1352_io_x2; // @[MUL.scala 102:19]
  wire  m_1352_io_x3; // @[MUL.scala 102:19]
  wire  m_1352_io_s; // @[MUL.scala 102:19]
  wire  m_1352_io_cout; // @[MUL.scala 102:19]
  wire  m_1353_io_x1; // @[MUL.scala 102:19]
  wire  m_1353_io_x2; // @[MUL.scala 102:19]
  wire  m_1353_io_x3; // @[MUL.scala 102:19]
  wire  m_1353_io_s; // @[MUL.scala 102:19]
  wire  m_1353_io_cout; // @[MUL.scala 102:19]
  wire  m_1354_io_x1; // @[MUL.scala 102:19]
  wire  m_1354_io_x2; // @[MUL.scala 102:19]
  wire  m_1354_io_x3; // @[MUL.scala 102:19]
  wire  m_1354_io_s; // @[MUL.scala 102:19]
  wire  m_1354_io_cout; // @[MUL.scala 102:19]
  wire  m_1355_io_x1; // @[MUL.scala 102:19]
  wire  m_1355_io_x2; // @[MUL.scala 102:19]
  wire  m_1355_io_x3; // @[MUL.scala 102:19]
  wire  m_1355_io_s; // @[MUL.scala 102:19]
  wire  m_1355_io_cout; // @[MUL.scala 102:19]
  wire  m_1356_io_x1; // @[MUL.scala 102:19]
  wire  m_1356_io_x2; // @[MUL.scala 102:19]
  wire  m_1356_io_x3; // @[MUL.scala 102:19]
  wire  m_1356_io_s; // @[MUL.scala 102:19]
  wire  m_1356_io_cout; // @[MUL.scala 102:19]
  wire  m_1357_io_x1; // @[MUL.scala 102:19]
  wire  m_1357_io_x2; // @[MUL.scala 102:19]
  wire  m_1357_io_x3; // @[MUL.scala 102:19]
  wire  m_1357_io_s; // @[MUL.scala 102:19]
  wire  m_1357_io_cout; // @[MUL.scala 102:19]
  wire  m_1358_io_x1; // @[MUL.scala 102:19]
  wire  m_1358_io_x2; // @[MUL.scala 102:19]
  wire  m_1358_io_x3; // @[MUL.scala 102:19]
  wire  m_1358_io_s; // @[MUL.scala 102:19]
  wire  m_1358_io_cout; // @[MUL.scala 102:19]
  wire  m_1359_io_x1; // @[MUL.scala 102:19]
  wire  m_1359_io_x2; // @[MUL.scala 102:19]
  wire  m_1359_io_x3; // @[MUL.scala 102:19]
  wire  m_1359_io_s; // @[MUL.scala 102:19]
  wire  m_1359_io_cout; // @[MUL.scala 102:19]
  wire  m_1360_io_x1; // @[MUL.scala 102:19]
  wire  m_1360_io_x2; // @[MUL.scala 102:19]
  wire  m_1360_io_x3; // @[MUL.scala 102:19]
  wire  m_1360_io_s; // @[MUL.scala 102:19]
  wire  m_1360_io_cout; // @[MUL.scala 102:19]
  wire  m_1361_io_x1; // @[MUL.scala 102:19]
  wire  m_1361_io_x2; // @[MUL.scala 102:19]
  wire  m_1361_io_x3; // @[MUL.scala 102:19]
  wire  m_1361_io_s; // @[MUL.scala 102:19]
  wire  m_1361_io_cout; // @[MUL.scala 102:19]
  wire  m_1362_io_x1; // @[MUL.scala 102:19]
  wire  m_1362_io_x2; // @[MUL.scala 102:19]
  wire  m_1362_io_x3; // @[MUL.scala 102:19]
  wire  m_1362_io_s; // @[MUL.scala 102:19]
  wire  m_1362_io_cout; // @[MUL.scala 102:19]
  wire  m_1363_io_x1; // @[MUL.scala 102:19]
  wire  m_1363_io_x2; // @[MUL.scala 102:19]
  wire  m_1363_io_x3; // @[MUL.scala 102:19]
  wire  m_1363_io_s; // @[MUL.scala 102:19]
  wire  m_1363_io_cout; // @[MUL.scala 102:19]
  wire  m_1364_io_x1; // @[MUL.scala 102:19]
  wire  m_1364_io_x2; // @[MUL.scala 102:19]
  wire  m_1364_io_x3; // @[MUL.scala 102:19]
  wire  m_1364_io_s; // @[MUL.scala 102:19]
  wire  m_1364_io_cout; // @[MUL.scala 102:19]
  wire  m_1365_io_x1; // @[MUL.scala 102:19]
  wire  m_1365_io_x2; // @[MUL.scala 102:19]
  wire  m_1365_io_x3; // @[MUL.scala 102:19]
  wire  m_1365_io_s; // @[MUL.scala 102:19]
  wire  m_1365_io_cout; // @[MUL.scala 102:19]
  wire  m_1366_io_x1; // @[MUL.scala 102:19]
  wire  m_1366_io_x2; // @[MUL.scala 102:19]
  wire  m_1366_io_x3; // @[MUL.scala 102:19]
  wire  m_1366_io_s; // @[MUL.scala 102:19]
  wire  m_1366_io_cout; // @[MUL.scala 102:19]
  wire  m_1367_io_x1; // @[MUL.scala 102:19]
  wire  m_1367_io_x2; // @[MUL.scala 102:19]
  wire  m_1367_io_x3; // @[MUL.scala 102:19]
  wire  m_1367_io_s; // @[MUL.scala 102:19]
  wire  m_1367_io_cout; // @[MUL.scala 102:19]
  wire  m_1368_io_x1; // @[MUL.scala 102:19]
  wire  m_1368_io_x2; // @[MUL.scala 102:19]
  wire  m_1368_io_x3; // @[MUL.scala 102:19]
  wire  m_1368_io_s; // @[MUL.scala 102:19]
  wire  m_1368_io_cout; // @[MUL.scala 102:19]
  wire  m_1369_io_x1; // @[MUL.scala 102:19]
  wire  m_1369_io_x2; // @[MUL.scala 102:19]
  wire  m_1369_io_x3; // @[MUL.scala 102:19]
  wire  m_1369_io_s; // @[MUL.scala 102:19]
  wire  m_1369_io_cout; // @[MUL.scala 102:19]
  wire  m_1370_io_x1; // @[MUL.scala 102:19]
  wire  m_1370_io_x2; // @[MUL.scala 102:19]
  wire  m_1370_io_x3; // @[MUL.scala 102:19]
  wire  m_1370_io_s; // @[MUL.scala 102:19]
  wire  m_1370_io_cout; // @[MUL.scala 102:19]
  wire  m_1371_io_in_0; // @[MUL.scala 124:19]
  wire  m_1371_io_in_1; // @[MUL.scala 124:19]
  wire  m_1371_io_out_0; // @[MUL.scala 124:19]
  wire  m_1371_io_out_1; // @[MUL.scala 124:19]
  wire  m_1372_io_x1; // @[MUL.scala 102:19]
  wire  m_1372_io_x2; // @[MUL.scala 102:19]
  wire  m_1372_io_x3; // @[MUL.scala 102:19]
  wire  m_1372_io_s; // @[MUL.scala 102:19]
  wire  m_1372_io_cout; // @[MUL.scala 102:19]
  wire  m_1373_io_x1; // @[MUL.scala 102:19]
  wire  m_1373_io_x2; // @[MUL.scala 102:19]
  wire  m_1373_io_x3; // @[MUL.scala 102:19]
  wire  m_1373_io_s; // @[MUL.scala 102:19]
  wire  m_1373_io_cout; // @[MUL.scala 102:19]
  wire  m_1374_io_in_0; // @[MUL.scala 124:19]
  wire  m_1374_io_in_1; // @[MUL.scala 124:19]
  wire  m_1374_io_out_0; // @[MUL.scala 124:19]
  wire  m_1374_io_out_1; // @[MUL.scala 124:19]
  wire  m_1375_io_x1; // @[MUL.scala 102:19]
  wire  m_1375_io_x2; // @[MUL.scala 102:19]
  wire  m_1375_io_x3; // @[MUL.scala 102:19]
  wire  m_1375_io_s; // @[MUL.scala 102:19]
  wire  m_1375_io_cout; // @[MUL.scala 102:19]
  wire  m_1376_io_x1; // @[MUL.scala 102:19]
  wire  m_1376_io_x2; // @[MUL.scala 102:19]
  wire  m_1376_io_x3; // @[MUL.scala 102:19]
  wire  m_1376_io_s; // @[MUL.scala 102:19]
  wire  m_1376_io_cout; // @[MUL.scala 102:19]
  wire  m_1377_io_in_0; // @[MUL.scala 124:19]
  wire  m_1377_io_in_1; // @[MUL.scala 124:19]
  wire  m_1377_io_out_0; // @[MUL.scala 124:19]
  wire  m_1377_io_out_1; // @[MUL.scala 124:19]
  wire  m_1378_io_x1; // @[MUL.scala 102:19]
  wire  m_1378_io_x2; // @[MUL.scala 102:19]
  wire  m_1378_io_x3; // @[MUL.scala 102:19]
  wire  m_1378_io_s; // @[MUL.scala 102:19]
  wire  m_1378_io_cout; // @[MUL.scala 102:19]
  wire  m_1379_io_x1; // @[MUL.scala 102:19]
  wire  m_1379_io_x2; // @[MUL.scala 102:19]
  wire  m_1379_io_x3; // @[MUL.scala 102:19]
  wire  m_1379_io_s; // @[MUL.scala 102:19]
  wire  m_1379_io_cout; // @[MUL.scala 102:19]
  wire  m_1380_io_in_0; // @[MUL.scala 124:19]
  wire  m_1380_io_in_1; // @[MUL.scala 124:19]
  wire  m_1380_io_out_0; // @[MUL.scala 124:19]
  wire  m_1380_io_out_1; // @[MUL.scala 124:19]
  wire  m_1381_io_x1; // @[MUL.scala 102:19]
  wire  m_1381_io_x2; // @[MUL.scala 102:19]
  wire  m_1381_io_x3; // @[MUL.scala 102:19]
  wire  m_1381_io_s; // @[MUL.scala 102:19]
  wire  m_1381_io_cout; // @[MUL.scala 102:19]
  wire  m_1382_io_x1; // @[MUL.scala 102:19]
  wire  m_1382_io_x2; // @[MUL.scala 102:19]
  wire  m_1382_io_x3; // @[MUL.scala 102:19]
  wire  m_1382_io_s; // @[MUL.scala 102:19]
  wire  m_1382_io_cout; // @[MUL.scala 102:19]
  wire  m_1383_io_in_0; // @[MUL.scala 124:19]
  wire  m_1383_io_in_1; // @[MUL.scala 124:19]
  wire  m_1383_io_out_0; // @[MUL.scala 124:19]
  wire  m_1383_io_out_1; // @[MUL.scala 124:19]
  wire  m_1384_io_x1; // @[MUL.scala 102:19]
  wire  m_1384_io_x2; // @[MUL.scala 102:19]
  wire  m_1384_io_x3; // @[MUL.scala 102:19]
  wire  m_1384_io_s; // @[MUL.scala 102:19]
  wire  m_1384_io_cout; // @[MUL.scala 102:19]
  wire  m_1385_io_x1; // @[MUL.scala 102:19]
  wire  m_1385_io_x2; // @[MUL.scala 102:19]
  wire  m_1385_io_x3; // @[MUL.scala 102:19]
  wire  m_1385_io_s; // @[MUL.scala 102:19]
  wire  m_1385_io_cout; // @[MUL.scala 102:19]
  wire  m_1386_io_x1; // @[MUL.scala 102:19]
  wire  m_1386_io_x2; // @[MUL.scala 102:19]
  wire  m_1386_io_x3; // @[MUL.scala 102:19]
  wire  m_1386_io_s; // @[MUL.scala 102:19]
  wire  m_1386_io_cout; // @[MUL.scala 102:19]
  wire  m_1387_io_x1; // @[MUL.scala 102:19]
  wire  m_1387_io_x2; // @[MUL.scala 102:19]
  wire  m_1387_io_x3; // @[MUL.scala 102:19]
  wire  m_1387_io_s; // @[MUL.scala 102:19]
  wire  m_1387_io_cout; // @[MUL.scala 102:19]
  wire  m_1388_io_x1; // @[MUL.scala 102:19]
  wire  m_1388_io_x2; // @[MUL.scala 102:19]
  wire  m_1388_io_x3; // @[MUL.scala 102:19]
  wire  m_1388_io_s; // @[MUL.scala 102:19]
  wire  m_1388_io_cout; // @[MUL.scala 102:19]
  wire  m_1389_io_x1; // @[MUL.scala 102:19]
  wire  m_1389_io_x2; // @[MUL.scala 102:19]
  wire  m_1389_io_x3; // @[MUL.scala 102:19]
  wire  m_1389_io_s; // @[MUL.scala 102:19]
  wire  m_1389_io_cout; // @[MUL.scala 102:19]
  wire  m_1390_io_x1; // @[MUL.scala 102:19]
  wire  m_1390_io_x2; // @[MUL.scala 102:19]
  wire  m_1390_io_x3; // @[MUL.scala 102:19]
  wire  m_1390_io_s; // @[MUL.scala 102:19]
  wire  m_1390_io_cout; // @[MUL.scala 102:19]
  wire  m_1391_io_x1; // @[MUL.scala 102:19]
  wire  m_1391_io_x2; // @[MUL.scala 102:19]
  wire  m_1391_io_x3; // @[MUL.scala 102:19]
  wire  m_1391_io_s; // @[MUL.scala 102:19]
  wire  m_1391_io_cout; // @[MUL.scala 102:19]
  wire  m_1392_io_x1; // @[MUL.scala 102:19]
  wire  m_1392_io_x2; // @[MUL.scala 102:19]
  wire  m_1392_io_x3; // @[MUL.scala 102:19]
  wire  m_1392_io_s; // @[MUL.scala 102:19]
  wire  m_1392_io_cout; // @[MUL.scala 102:19]
  wire  m_1393_io_x1; // @[MUL.scala 102:19]
  wire  m_1393_io_x2; // @[MUL.scala 102:19]
  wire  m_1393_io_x3; // @[MUL.scala 102:19]
  wire  m_1393_io_s; // @[MUL.scala 102:19]
  wire  m_1393_io_cout; // @[MUL.scala 102:19]
  wire  m_1394_io_x1; // @[MUL.scala 102:19]
  wire  m_1394_io_x2; // @[MUL.scala 102:19]
  wire  m_1394_io_x3; // @[MUL.scala 102:19]
  wire  m_1394_io_s; // @[MUL.scala 102:19]
  wire  m_1394_io_cout; // @[MUL.scala 102:19]
  wire  m_1395_io_x1; // @[MUL.scala 102:19]
  wire  m_1395_io_x2; // @[MUL.scala 102:19]
  wire  m_1395_io_x3; // @[MUL.scala 102:19]
  wire  m_1395_io_s; // @[MUL.scala 102:19]
  wire  m_1395_io_cout; // @[MUL.scala 102:19]
  wire  m_1396_io_x1; // @[MUL.scala 102:19]
  wire  m_1396_io_x2; // @[MUL.scala 102:19]
  wire  m_1396_io_x3; // @[MUL.scala 102:19]
  wire  m_1396_io_s; // @[MUL.scala 102:19]
  wire  m_1396_io_cout; // @[MUL.scala 102:19]
  wire  m_1397_io_x1; // @[MUL.scala 102:19]
  wire  m_1397_io_x2; // @[MUL.scala 102:19]
  wire  m_1397_io_x3; // @[MUL.scala 102:19]
  wire  m_1397_io_s; // @[MUL.scala 102:19]
  wire  m_1397_io_cout; // @[MUL.scala 102:19]
  wire  m_1398_io_x1; // @[MUL.scala 102:19]
  wire  m_1398_io_x2; // @[MUL.scala 102:19]
  wire  m_1398_io_x3; // @[MUL.scala 102:19]
  wire  m_1398_io_s; // @[MUL.scala 102:19]
  wire  m_1398_io_cout; // @[MUL.scala 102:19]
  wire  m_1399_io_x1; // @[MUL.scala 102:19]
  wire  m_1399_io_x2; // @[MUL.scala 102:19]
  wire  m_1399_io_x3; // @[MUL.scala 102:19]
  wire  m_1399_io_s; // @[MUL.scala 102:19]
  wire  m_1399_io_cout; // @[MUL.scala 102:19]
  wire  m_1400_io_x1; // @[MUL.scala 102:19]
  wire  m_1400_io_x2; // @[MUL.scala 102:19]
  wire  m_1400_io_x3; // @[MUL.scala 102:19]
  wire  m_1400_io_s; // @[MUL.scala 102:19]
  wire  m_1400_io_cout; // @[MUL.scala 102:19]
  wire  m_1401_io_x1; // @[MUL.scala 102:19]
  wire  m_1401_io_x2; // @[MUL.scala 102:19]
  wire  m_1401_io_x3; // @[MUL.scala 102:19]
  wire  m_1401_io_s; // @[MUL.scala 102:19]
  wire  m_1401_io_cout; // @[MUL.scala 102:19]
  wire  m_1402_io_x1; // @[MUL.scala 102:19]
  wire  m_1402_io_x2; // @[MUL.scala 102:19]
  wire  m_1402_io_x3; // @[MUL.scala 102:19]
  wire  m_1402_io_s; // @[MUL.scala 102:19]
  wire  m_1402_io_cout; // @[MUL.scala 102:19]
  wire  m_1403_io_x1; // @[MUL.scala 102:19]
  wire  m_1403_io_x2; // @[MUL.scala 102:19]
  wire  m_1403_io_x3; // @[MUL.scala 102:19]
  wire  m_1403_io_s; // @[MUL.scala 102:19]
  wire  m_1403_io_cout; // @[MUL.scala 102:19]
  wire  m_1404_io_x1; // @[MUL.scala 102:19]
  wire  m_1404_io_x2; // @[MUL.scala 102:19]
  wire  m_1404_io_x3; // @[MUL.scala 102:19]
  wire  m_1404_io_s; // @[MUL.scala 102:19]
  wire  m_1404_io_cout; // @[MUL.scala 102:19]
  wire  m_1405_io_x1; // @[MUL.scala 102:19]
  wire  m_1405_io_x2; // @[MUL.scala 102:19]
  wire  m_1405_io_x3; // @[MUL.scala 102:19]
  wire  m_1405_io_s; // @[MUL.scala 102:19]
  wire  m_1405_io_cout; // @[MUL.scala 102:19]
  wire  m_1406_io_x1; // @[MUL.scala 102:19]
  wire  m_1406_io_x2; // @[MUL.scala 102:19]
  wire  m_1406_io_x3; // @[MUL.scala 102:19]
  wire  m_1406_io_s; // @[MUL.scala 102:19]
  wire  m_1406_io_cout; // @[MUL.scala 102:19]
  wire  m_1407_io_x1; // @[MUL.scala 102:19]
  wire  m_1407_io_x2; // @[MUL.scala 102:19]
  wire  m_1407_io_x3; // @[MUL.scala 102:19]
  wire  m_1407_io_s; // @[MUL.scala 102:19]
  wire  m_1407_io_cout; // @[MUL.scala 102:19]
  wire  m_1408_io_x1; // @[MUL.scala 102:19]
  wire  m_1408_io_x2; // @[MUL.scala 102:19]
  wire  m_1408_io_x3; // @[MUL.scala 102:19]
  wire  m_1408_io_s; // @[MUL.scala 102:19]
  wire  m_1408_io_cout; // @[MUL.scala 102:19]
  wire  m_1409_io_x1; // @[MUL.scala 102:19]
  wire  m_1409_io_x2; // @[MUL.scala 102:19]
  wire  m_1409_io_x3; // @[MUL.scala 102:19]
  wire  m_1409_io_s; // @[MUL.scala 102:19]
  wire  m_1409_io_cout; // @[MUL.scala 102:19]
  wire  m_1410_io_x1; // @[MUL.scala 102:19]
  wire  m_1410_io_x2; // @[MUL.scala 102:19]
  wire  m_1410_io_x3; // @[MUL.scala 102:19]
  wire  m_1410_io_s; // @[MUL.scala 102:19]
  wire  m_1410_io_cout; // @[MUL.scala 102:19]
  wire  m_1411_io_x1; // @[MUL.scala 102:19]
  wire  m_1411_io_x2; // @[MUL.scala 102:19]
  wire  m_1411_io_x3; // @[MUL.scala 102:19]
  wire  m_1411_io_s; // @[MUL.scala 102:19]
  wire  m_1411_io_cout; // @[MUL.scala 102:19]
  wire  m_1412_io_x1; // @[MUL.scala 102:19]
  wire  m_1412_io_x2; // @[MUL.scala 102:19]
  wire  m_1412_io_x3; // @[MUL.scala 102:19]
  wire  m_1412_io_s; // @[MUL.scala 102:19]
  wire  m_1412_io_cout; // @[MUL.scala 102:19]
  wire  m_1413_io_x1; // @[MUL.scala 102:19]
  wire  m_1413_io_x2; // @[MUL.scala 102:19]
  wire  m_1413_io_x3; // @[MUL.scala 102:19]
  wire  m_1413_io_s; // @[MUL.scala 102:19]
  wire  m_1413_io_cout; // @[MUL.scala 102:19]
  wire  m_1414_io_in_0; // @[MUL.scala 124:19]
  wire  m_1414_io_in_1; // @[MUL.scala 124:19]
  wire  m_1414_io_out_0; // @[MUL.scala 124:19]
  wire  m_1414_io_out_1; // @[MUL.scala 124:19]
  wire  m_1415_io_x1; // @[MUL.scala 102:19]
  wire  m_1415_io_x2; // @[MUL.scala 102:19]
  wire  m_1415_io_x3; // @[MUL.scala 102:19]
  wire  m_1415_io_s; // @[MUL.scala 102:19]
  wire  m_1415_io_cout; // @[MUL.scala 102:19]
  wire  m_1416_io_x1; // @[MUL.scala 102:19]
  wire  m_1416_io_x2; // @[MUL.scala 102:19]
  wire  m_1416_io_x3; // @[MUL.scala 102:19]
  wire  m_1416_io_s; // @[MUL.scala 102:19]
  wire  m_1416_io_cout; // @[MUL.scala 102:19]
  wire  m_1417_io_x1; // @[MUL.scala 102:19]
  wire  m_1417_io_x2; // @[MUL.scala 102:19]
  wire  m_1417_io_x3; // @[MUL.scala 102:19]
  wire  m_1417_io_s; // @[MUL.scala 102:19]
  wire  m_1417_io_cout; // @[MUL.scala 102:19]
  wire  m_1418_io_in_0; // @[MUL.scala 124:19]
  wire  m_1418_io_in_1; // @[MUL.scala 124:19]
  wire  m_1418_io_out_0; // @[MUL.scala 124:19]
  wire  m_1418_io_out_1; // @[MUL.scala 124:19]
  wire  m_1419_io_x1; // @[MUL.scala 102:19]
  wire  m_1419_io_x2; // @[MUL.scala 102:19]
  wire  m_1419_io_x3; // @[MUL.scala 102:19]
  wire  m_1419_io_s; // @[MUL.scala 102:19]
  wire  m_1419_io_cout; // @[MUL.scala 102:19]
  wire  m_1420_io_x1; // @[MUL.scala 102:19]
  wire  m_1420_io_x2; // @[MUL.scala 102:19]
  wire  m_1420_io_x3; // @[MUL.scala 102:19]
  wire  m_1420_io_s; // @[MUL.scala 102:19]
  wire  m_1420_io_cout; // @[MUL.scala 102:19]
  wire  m_1421_io_x1; // @[MUL.scala 102:19]
  wire  m_1421_io_x2; // @[MUL.scala 102:19]
  wire  m_1421_io_x3; // @[MUL.scala 102:19]
  wire  m_1421_io_s; // @[MUL.scala 102:19]
  wire  m_1421_io_cout; // @[MUL.scala 102:19]
  wire  m_1422_io_in_0; // @[MUL.scala 124:19]
  wire  m_1422_io_in_1; // @[MUL.scala 124:19]
  wire  m_1422_io_out_0; // @[MUL.scala 124:19]
  wire  m_1422_io_out_1; // @[MUL.scala 124:19]
  wire  m_1423_io_x1; // @[MUL.scala 102:19]
  wire  m_1423_io_x2; // @[MUL.scala 102:19]
  wire  m_1423_io_x3; // @[MUL.scala 102:19]
  wire  m_1423_io_s; // @[MUL.scala 102:19]
  wire  m_1423_io_cout; // @[MUL.scala 102:19]
  wire  m_1424_io_x1; // @[MUL.scala 102:19]
  wire  m_1424_io_x2; // @[MUL.scala 102:19]
  wire  m_1424_io_x3; // @[MUL.scala 102:19]
  wire  m_1424_io_s; // @[MUL.scala 102:19]
  wire  m_1424_io_cout; // @[MUL.scala 102:19]
  wire  m_1425_io_x1; // @[MUL.scala 102:19]
  wire  m_1425_io_x2; // @[MUL.scala 102:19]
  wire  m_1425_io_x3; // @[MUL.scala 102:19]
  wire  m_1425_io_s; // @[MUL.scala 102:19]
  wire  m_1425_io_cout; // @[MUL.scala 102:19]
  wire  m_1426_io_in_0; // @[MUL.scala 124:19]
  wire  m_1426_io_in_1; // @[MUL.scala 124:19]
  wire  m_1426_io_out_0; // @[MUL.scala 124:19]
  wire  m_1426_io_out_1; // @[MUL.scala 124:19]
  wire  m_1427_io_x1; // @[MUL.scala 102:19]
  wire  m_1427_io_x2; // @[MUL.scala 102:19]
  wire  m_1427_io_x3; // @[MUL.scala 102:19]
  wire  m_1427_io_s; // @[MUL.scala 102:19]
  wire  m_1427_io_cout; // @[MUL.scala 102:19]
  wire  m_1428_io_x1; // @[MUL.scala 102:19]
  wire  m_1428_io_x2; // @[MUL.scala 102:19]
  wire  m_1428_io_x3; // @[MUL.scala 102:19]
  wire  m_1428_io_s; // @[MUL.scala 102:19]
  wire  m_1428_io_cout; // @[MUL.scala 102:19]
  wire  m_1429_io_x1; // @[MUL.scala 102:19]
  wire  m_1429_io_x2; // @[MUL.scala 102:19]
  wire  m_1429_io_x3; // @[MUL.scala 102:19]
  wire  m_1429_io_s; // @[MUL.scala 102:19]
  wire  m_1429_io_cout; // @[MUL.scala 102:19]
  wire  m_1430_io_x1; // @[MUL.scala 102:19]
  wire  m_1430_io_x2; // @[MUL.scala 102:19]
  wire  m_1430_io_x3; // @[MUL.scala 102:19]
  wire  m_1430_io_s; // @[MUL.scala 102:19]
  wire  m_1430_io_cout; // @[MUL.scala 102:19]
  wire  m_1431_io_x1; // @[MUL.scala 102:19]
  wire  m_1431_io_x2; // @[MUL.scala 102:19]
  wire  m_1431_io_x3; // @[MUL.scala 102:19]
  wire  m_1431_io_s; // @[MUL.scala 102:19]
  wire  m_1431_io_cout; // @[MUL.scala 102:19]
  wire  m_1432_io_x1; // @[MUL.scala 102:19]
  wire  m_1432_io_x2; // @[MUL.scala 102:19]
  wire  m_1432_io_x3; // @[MUL.scala 102:19]
  wire  m_1432_io_s; // @[MUL.scala 102:19]
  wire  m_1432_io_cout; // @[MUL.scala 102:19]
  wire  m_1433_io_x1; // @[MUL.scala 102:19]
  wire  m_1433_io_x2; // @[MUL.scala 102:19]
  wire  m_1433_io_x3; // @[MUL.scala 102:19]
  wire  m_1433_io_s; // @[MUL.scala 102:19]
  wire  m_1433_io_cout; // @[MUL.scala 102:19]
  wire  m_1434_io_x1; // @[MUL.scala 102:19]
  wire  m_1434_io_x2; // @[MUL.scala 102:19]
  wire  m_1434_io_x3; // @[MUL.scala 102:19]
  wire  m_1434_io_s; // @[MUL.scala 102:19]
  wire  m_1434_io_cout; // @[MUL.scala 102:19]
  wire  m_1435_io_x1; // @[MUL.scala 102:19]
  wire  m_1435_io_x2; // @[MUL.scala 102:19]
  wire  m_1435_io_x3; // @[MUL.scala 102:19]
  wire  m_1435_io_s; // @[MUL.scala 102:19]
  wire  m_1435_io_cout; // @[MUL.scala 102:19]
  wire  m_1436_io_x1; // @[MUL.scala 102:19]
  wire  m_1436_io_x2; // @[MUL.scala 102:19]
  wire  m_1436_io_x3; // @[MUL.scala 102:19]
  wire  m_1436_io_s; // @[MUL.scala 102:19]
  wire  m_1436_io_cout; // @[MUL.scala 102:19]
  wire  m_1437_io_x1; // @[MUL.scala 102:19]
  wire  m_1437_io_x2; // @[MUL.scala 102:19]
  wire  m_1437_io_x3; // @[MUL.scala 102:19]
  wire  m_1437_io_s; // @[MUL.scala 102:19]
  wire  m_1437_io_cout; // @[MUL.scala 102:19]
  wire  m_1438_io_x1; // @[MUL.scala 102:19]
  wire  m_1438_io_x2; // @[MUL.scala 102:19]
  wire  m_1438_io_x3; // @[MUL.scala 102:19]
  wire  m_1438_io_s; // @[MUL.scala 102:19]
  wire  m_1438_io_cout; // @[MUL.scala 102:19]
  wire  m_1439_io_x1; // @[MUL.scala 102:19]
  wire  m_1439_io_x2; // @[MUL.scala 102:19]
  wire  m_1439_io_x3; // @[MUL.scala 102:19]
  wire  m_1439_io_s; // @[MUL.scala 102:19]
  wire  m_1439_io_cout; // @[MUL.scala 102:19]
  wire  m_1440_io_x1; // @[MUL.scala 102:19]
  wire  m_1440_io_x2; // @[MUL.scala 102:19]
  wire  m_1440_io_x3; // @[MUL.scala 102:19]
  wire  m_1440_io_s; // @[MUL.scala 102:19]
  wire  m_1440_io_cout; // @[MUL.scala 102:19]
  wire  m_1441_io_x1; // @[MUL.scala 102:19]
  wire  m_1441_io_x2; // @[MUL.scala 102:19]
  wire  m_1441_io_x3; // @[MUL.scala 102:19]
  wire  m_1441_io_s; // @[MUL.scala 102:19]
  wire  m_1441_io_cout; // @[MUL.scala 102:19]
  wire  m_1442_io_x1; // @[MUL.scala 102:19]
  wire  m_1442_io_x2; // @[MUL.scala 102:19]
  wire  m_1442_io_x3; // @[MUL.scala 102:19]
  wire  m_1442_io_s; // @[MUL.scala 102:19]
  wire  m_1442_io_cout; // @[MUL.scala 102:19]
  wire  m_1443_io_x1; // @[MUL.scala 102:19]
  wire  m_1443_io_x2; // @[MUL.scala 102:19]
  wire  m_1443_io_x3; // @[MUL.scala 102:19]
  wire  m_1443_io_s; // @[MUL.scala 102:19]
  wire  m_1443_io_cout; // @[MUL.scala 102:19]
  wire  m_1444_io_x1; // @[MUL.scala 102:19]
  wire  m_1444_io_x2; // @[MUL.scala 102:19]
  wire  m_1444_io_x3; // @[MUL.scala 102:19]
  wire  m_1444_io_s; // @[MUL.scala 102:19]
  wire  m_1444_io_cout; // @[MUL.scala 102:19]
  wire  m_1445_io_x1; // @[MUL.scala 102:19]
  wire  m_1445_io_x2; // @[MUL.scala 102:19]
  wire  m_1445_io_x3; // @[MUL.scala 102:19]
  wire  m_1445_io_s; // @[MUL.scala 102:19]
  wire  m_1445_io_cout; // @[MUL.scala 102:19]
  wire  m_1446_io_x1; // @[MUL.scala 102:19]
  wire  m_1446_io_x2; // @[MUL.scala 102:19]
  wire  m_1446_io_x3; // @[MUL.scala 102:19]
  wire  m_1446_io_s; // @[MUL.scala 102:19]
  wire  m_1446_io_cout; // @[MUL.scala 102:19]
  wire  m_1447_io_x1; // @[MUL.scala 102:19]
  wire  m_1447_io_x2; // @[MUL.scala 102:19]
  wire  m_1447_io_x3; // @[MUL.scala 102:19]
  wire  m_1447_io_s; // @[MUL.scala 102:19]
  wire  m_1447_io_cout; // @[MUL.scala 102:19]
  wire  m_1448_io_x1; // @[MUL.scala 102:19]
  wire  m_1448_io_x2; // @[MUL.scala 102:19]
  wire  m_1448_io_x3; // @[MUL.scala 102:19]
  wire  m_1448_io_s; // @[MUL.scala 102:19]
  wire  m_1448_io_cout; // @[MUL.scala 102:19]
  wire  m_1449_io_x1; // @[MUL.scala 102:19]
  wire  m_1449_io_x2; // @[MUL.scala 102:19]
  wire  m_1449_io_x3; // @[MUL.scala 102:19]
  wire  m_1449_io_s; // @[MUL.scala 102:19]
  wire  m_1449_io_cout; // @[MUL.scala 102:19]
  wire  m_1450_io_x1; // @[MUL.scala 102:19]
  wire  m_1450_io_x2; // @[MUL.scala 102:19]
  wire  m_1450_io_x3; // @[MUL.scala 102:19]
  wire  m_1450_io_s; // @[MUL.scala 102:19]
  wire  m_1450_io_cout; // @[MUL.scala 102:19]
  wire  m_1451_io_x1; // @[MUL.scala 102:19]
  wire  m_1451_io_x2; // @[MUL.scala 102:19]
  wire  m_1451_io_x3; // @[MUL.scala 102:19]
  wire  m_1451_io_s; // @[MUL.scala 102:19]
  wire  m_1451_io_cout; // @[MUL.scala 102:19]
  wire  m_1452_io_x1; // @[MUL.scala 102:19]
  wire  m_1452_io_x2; // @[MUL.scala 102:19]
  wire  m_1452_io_x3; // @[MUL.scala 102:19]
  wire  m_1452_io_s; // @[MUL.scala 102:19]
  wire  m_1452_io_cout; // @[MUL.scala 102:19]
  wire  m_1453_io_x1; // @[MUL.scala 102:19]
  wire  m_1453_io_x2; // @[MUL.scala 102:19]
  wire  m_1453_io_x3; // @[MUL.scala 102:19]
  wire  m_1453_io_s; // @[MUL.scala 102:19]
  wire  m_1453_io_cout; // @[MUL.scala 102:19]
  wire  m_1454_io_x1; // @[MUL.scala 102:19]
  wire  m_1454_io_x2; // @[MUL.scala 102:19]
  wire  m_1454_io_x3; // @[MUL.scala 102:19]
  wire  m_1454_io_s; // @[MUL.scala 102:19]
  wire  m_1454_io_cout; // @[MUL.scala 102:19]
  wire  m_1455_io_x1; // @[MUL.scala 102:19]
  wire  m_1455_io_x2; // @[MUL.scala 102:19]
  wire  m_1455_io_x3; // @[MUL.scala 102:19]
  wire  m_1455_io_s; // @[MUL.scala 102:19]
  wire  m_1455_io_cout; // @[MUL.scala 102:19]
  wire  m_1456_io_x1; // @[MUL.scala 102:19]
  wire  m_1456_io_x2; // @[MUL.scala 102:19]
  wire  m_1456_io_x3; // @[MUL.scala 102:19]
  wire  m_1456_io_s; // @[MUL.scala 102:19]
  wire  m_1456_io_cout; // @[MUL.scala 102:19]
  wire  m_1457_io_x1; // @[MUL.scala 102:19]
  wire  m_1457_io_x2; // @[MUL.scala 102:19]
  wire  m_1457_io_x3; // @[MUL.scala 102:19]
  wire  m_1457_io_s; // @[MUL.scala 102:19]
  wire  m_1457_io_cout; // @[MUL.scala 102:19]
  wire  m_1458_io_x1; // @[MUL.scala 102:19]
  wire  m_1458_io_x2; // @[MUL.scala 102:19]
  wire  m_1458_io_x3; // @[MUL.scala 102:19]
  wire  m_1458_io_s; // @[MUL.scala 102:19]
  wire  m_1458_io_cout; // @[MUL.scala 102:19]
  wire  m_1459_io_x1; // @[MUL.scala 102:19]
  wire  m_1459_io_x2; // @[MUL.scala 102:19]
  wire  m_1459_io_x3; // @[MUL.scala 102:19]
  wire  m_1459_io_s; // @[MUL.scala 102:19]
  wire  m_1459_io_cout; // @[MUL.scala 102:19]
  wire  m_1460_io_x1; // @[MUL.scala 102:19]
  wire  m_1460_io_x2; // @[MUL.scala 102:19]
  wire  m_1460_io_x3; // @[MUL.scala 102:19]
  wire  m_1460_io_s; // @[MUL.scala 102:19]
  wire  m_1460_io_cout; // @[MUL.scala 102:19]
  wire  m_1461_io_x1; // @[MUL.scala 102:19]
  wire  m_1461_io_x2; // @[MUL.scala 102:19]
  wire  m_1461_io_x3; // @[MUL.scala 102:19]
  wire  m_1461_io_s; // @[MUL.scala 102:19]
  wire  m_1461_io_cout; // @[MUL.scala 102:19]
  wire  m_1462_io_x1; // @[MUL.scala 102:19]
  wire  m_1462_io_x2; // @[MUL.scala 102:19]
  wire  m_1462_io_x3; // @[MUL.scala 102:19]
  wire  m_1462_io_s; // @[MUL.scala 102:19]
  wire  m_1462_io_cout; // @[MUL.scala 102:19]
  wire  m_1463_io_x1; // @[MUL.scala 102:19]
  wire  m_1463_io_x2; // @[MUL.scala 102:19]
  wire  m_1463_io_x3; // @[MUL.scala 102:19]
  wire  m_1463_io_s; // @[MUL.scala 102:19]
  wire  m_1463_io_cout; // @[MUL.scala 102:19]
  wire  m_1464_io_x1; // @[MUL.scala 102:19]
  wire  m_1464_io_x2; // @[MUL.scala 102:19]
  wire  m_1464_io_x3; // @[MUL.scala 102:19]
  wire  m_1464_io_s; // @[MUL.scala 102:19]
  wire  m_1464_io_cout; // @[MUL.scala 102:19]
  wire  m_1465_io_x1; // @[MUL.scala 102:19]
  wire  m_1465_io_x2; // @[MUL.scala 102:19]
  wire  m_1465_io_x3; // @[MUL.scala 102:19]
  wire  m_1465_io_s; // @[MUL.scala 102:19]
  wire  m_1465_io_cout; // @[MUL.scala 102:19]
  wire  m_1466_io_x1; // @[MUL.scala 102:19]
  wire  m_1466_io_x2; // @[MUL.scala 102:19]
  wire  m_1466_io_x3; // @[MUL.scala 102:19]
  wire  m_1466_io_s; // @[MUL.scala 102:19]
  wire  m_1466_io_cout; // @[MUL.scala 102:19]
  wire  m_1467_io_in_0; // @[MUL.scala 124:19]
  wire  m_1467_io_in_1; // @[MUL.scala 124:19]
  wire  m_1467_io_out_0; // @[MUL.scala 124:19]
  wire  m_1467_io_out_1; // @[MUL.scala 124:19]
  wire  m_1468_io_x1; // @[MUL.scala 102:19]
  wire  m_1468_io_x2; // @[MUL.scala 102:19]
  wire  m_1468_io_x3; // @[MUL.scala 102:19]
  wire  m_1468_io_s; // @[MUL.scala 102:19]
  wire  m_1468_io_cout; // @[MUL.scala 102:19]
  wire  m_1469_io_x1; // @[MUL.scala 102:19]
  wire  m_1469_io_x2; // @[MUL.scala 102:19]
  wire  m_1469_io_x3; // @[MUL.scala 102:19]
  wire  m_1469_io_s; // @[MUL.scala 102:19]
  wire  m_1469_io_cout; // @[MUL.scala 102:19]
  wire  m_1470_io_x1; // @[MUL.scala 102:19]
  wire  m_1470_io_x2; // @[MUL.scala 102:19]
  wire  m_1470_io_x3; // @[MUL.scala 102:19]
  wire  m_1470_io_s; // @[MUL.scala 102:19]
  wire  m_1470_io_cout; // @[MUL.scala 102:19]
  wire  m_1471_io_x1; // @[MUL.scala 102:19]
  wire  m_1471_io_x2; // @[MUL.scala 102:19]
  wire  m_1471_io_x3; // @[MUL.scala 102:19]
  wire  m_1471_io_s; // @[MUL.scala 102:19]
  wire  m_1471_io_cout; // @[MUL.scala 102:19]
  wire  m_1472_io_in_0; // @[MUL.scala 124:19]
  wire  m_1472_io_in_1; // @[MUL.scala 124:19]
  wire  m_1472_io_out_0; // @[MUL.scala 124:19]
  wire  m_1472_io_out_1; // @[MUL.scala 124:19]
  wire  m_1473_io_x1; // @[MUL.scala 102:19]
  wire  m_1473_io_x2; // @[MUL.scala 102:19]
  wire  m_1473_io_x3; // @[MUL.scala 102:19]
  wire  m_1473_io_s; // @[MUL.scala 102:19]
  wire  m_1473_io_cout; // @[MUL.scala 102:19]
  wire  m_1474_io_x1; // @[MUL.scala 102:19]
  wire  m_1474_io_x2; // @[MUL.scala 102:19]
  wire  m_1474_io_x3; // @[MUL.scala 102:19]
  wire  m_1474_io_s; // @[MUL.scala 102:19]
  wire  m_1474_io_cout; // @[MUL.scala 102:19]
  wire  m_1475_io_x1; // @[MUL.scala 102:19]
  wire  m_1475_io_x2; // @[MUL.scala 102:19]
  wire  m_1475_io_x3; // @[MUL.scala 102:19]
  wire  m_1475_io_s; // @[MUL.scala 102:19]
  wire  m_1475_io_cout; // @[MUL.scala 102:19]
  wire  m_1476_io_x1; // @[MUL.scala 102:19]
  wire  m_1476_io_x2; // @[MUL.scala 102:19]
  wire  m_1476_io_x3; // @[MUL.scala 102:19]
  wire  m_1476_io_s; // @[MUL.scala 102:19]
  wire  m_1476_io_cout; // @[MUL.scala 102:19]
  wire  m_1477_io_in_0; // @[MUL.scala 124:19]
  wire  m_1477_io_in_1; // @[MUL.scala 124:19]
  wire  m_1477_io_out_0; // @[MUL.scala 124:19]
  wire  m_1477_io_out_1; // @[MUL.scala 124:19]
  wire  m_1478_io_x1; // @[MUL.scala 102:19]
  wire  m_1478_io_x2; // @[MUL.scala 102:19]
  wire  m_1478_io_x3; // @[MUL.scala 102:19]
  wire  m_1478_io_s; // @[MUL.scala 102:19]
  wire  m_1478_io_cout; // @[MUL.scala 102:19]
  wire  m_1479_io_x1; // @[MUL.scala 102:19]
  wire  m_1479_io_x2; // @[MUL.scala 102:19]
  wire  m_1479_io_x3; // @[MUL.scala 102:19]
  wire  m_1479_io_s; // @[MUL.scala 102:19]
  wire  m_1479_io_cout; // @[MUL.scala 102:19]
  wire  m_1480_io_x1; // @[MUL.scala 102:19]
  wire  m_1480_io_x2; // @[MUL.scala 102:19]
  wire  m_1480_io_x3; // @[MUL.scala 102:19]
  wire  m_1480_io_s; // @[MUL.scala 102:19]
  wire  m_1480_io_cout; // @[MUL.scala 102:19]
  wire  m_1481_io_x1; // @[MUL.scala 102:19]
  wire  m_1481_io_x2; // @[MUL.scala 102:19]
  wire  m_1481_io_x3; // @[MUL.scala 102:19]
  wire  m_1481_io_s; // @[MUL.scala 102:19]
  wire  m_1481_io_cout; // @[MUL.scala 102:19]
  wire  m_1482_io_in_0; // @[MUL.scala 124:19]
  wire  m_1482_io_in_1; // @[MUL.scala 124:19]
  wire  m_1482_io_out_0; // @[MUL.scala 124:19]
  wire  m_1482_io_out_1; // @[MUL.scala 124:19]
  wire  m_1483_io_x1; // @[MUL.scala 102:19]
  wire  m_1483_io_x2; // @[MUL.scala 102:19]
  wire  m_1483_io_x3; // @[MUL.scala 102:19]
  wire  m_1483_io_s; // @[MUL.scala 102:19]
  wire  m_1483_io_cout; // @[MUL.scala 102:19]
  wire  m_1484_io_x1; // @[MUL.scala 102:19]
  wire  m_1484_io_x2; // @[MUL.scala 102:19]
  wire  m_1484_io_x3; // @[MUL.scala 102:19]
  wire  m_1484_io_s; // @[MUL.scala 102:19]
  wire  m_1484_io_cout; // @[MUL.scala 102:19]
  wire  m_1485_io_x1; // @[MUL.scala 102:19]
  wire  m_1485_io_x2; // @[MUL.scala 102:19]
  wire  m_1485_io_x3; // @[MUL.scala 102:19]
  wire  m_1485_io_s; // @[MUL.scala 102:19]
  wire  m_1485_io_cout; // @[MUL.scala 102:19]
  wire  m_1486_io_x1; // @[MUL.scala 102:19]
  wire  m_1486_io_x2; // @[MUL.scala 102:19]
  wire  m_1486_io_x3; // @[MUL.scala 102:19]
  wire  m_1486_io_s; // @[MUL.scala 102:19]
  wire  m_1486_io_cout; // @[MUL.scala 102:19]
  wire  m_1487_io_in_0; // @[MUL.scala 124:19]
  wire  m_1487_io_in_1; // @[MUL.scala 124:19]
  wire  m_1487_io_out_0; // @[MUL.scala 124:19]
  wire  m_1487_io_out_1; // @[MUL.scala 124:19]
  wire  m_1488_io_x1; // @[MUL.scala 102:19]
  wire  m_1488_io_x2; // @[MUL.scala 102:19]
  wire  m_1488_io_x3; // @[MUL.scala 102:19]
  wire  m_1488_io_s; // @[MUL.scala 102:19]
  wire  m_1488_io_cout; // @[MUL.scala 102:19]
  wire  m_1489_io_x1; // @[MUL.scala 102:19]
  wire  m_1489_io_x2; // @[MUL.scala 102:19]
  wire  m_1489_io_x3; // @[MUL.scala 102:19]
  wire  m_1489_io_s; // @[MUL.scala 102:19]
  wire  m_1489_io_cout; // @[MUL.scala 102:19]
  wire  m_1490_io_x1; // @[MUL.scala 102:19]
  wire  m_1490_io_x2; // @[MUL.scala 102:19]
  wire  m_1490_io_x3; // @[MUL.scala 102:19]
  wire  m_1490_io_s; // @[MUL.scala 102:19]
  wire  m_1490_io_cout; // @[MUL.scala 102:19]
  wire  m_1491_io_x1; // @[MUL.scala 102:19]
  wire  m_1491_io_x2; // @[MUL.scala 102:19]
  wire  m_1491_io_x3; // @[MUL.scala 102:19]
  wire  m_1491_io_s; // @[MUL.scala 102:19]
  wire  m_1491_io_cout; // @[MUL.scala 102:19]
  wire  m_1492_io_x1; // @[MUL.scala 102:19]
  wire  m_1492_io_x2; // @[MUL.scala 102:19]
  wire  m_1492_io_x3; // @[MUL.scala 102:19]
  wire  m_1492_io_s; // @[MUL.scala 102:19]
  wire  m_1492_io_cout; // @[MUL.scala 102:19]
  wire  m_1493_io_x1; // @[MUL.scala 102:19]
  wire  m_1493_io_x2; // @[MUL.scala 102:19]
  wire  m_1493_io_x3; // @[MUL.scala 102:19]
  wire  m_1493_io_s; // @[MUL.scala 102:19]
  wire  m_1493_io_cout; // @[MUL.scala 102:19]
  wire  m_1494_io_x1; // @[MUL.scala 102:19]
  wire  m_1494_io_x2; // @[MUL.scala 102:19]
  wire  m_1494_io_x3; // @[MUL.scala 102:19]
  wire  m_1494_io_s; // @[MUL.scala 102:19]
  wire  m_1494_io_cout; // @[MUL.scala 102:19]
  wire  m_1495_io_x1; // @[MUL.scala 102:19]
  wire  m_1495_io_x2; // @[MUL.scala 102:19]
  wire  m_1495_io_x3; // @[MUL.scala 102:19]
  wire  m_1495_io_s; // @[MUL.scala 102:19]
  wire  m_1495_io_cout; // @[MUL.scala 102:19]
  wire  m_1496_io_x1; // @[MUL.scala 102:19]
  wire  m_1496_io_x2; // @[MUL.scala 102:19]
  wire  m_1496_io_x3; // @[MUL.scala 102:19]
  wire  m_1496_io_s; // @[MUL.scala 102:19]
  wire  m_1496_io_cout; // @[MUL.scala 102:19]
  wire  m_1497_io_x1; // @[MUL.scala 102:19]
  wire  m_1497_io_x2; // @[MUL.scala 102:19]
  wire  m_1497_io_x3; // @[MUL.scala 102:19]
  wire  m_1497_io_s; // @[MUL.scala 102:19]
  wire  m_1497_io_cout; // @[MUL.scala 102:19]
  wire  m_1498_io_x1; // @[MUL.scala 102:19]
  wire  m_1498_io_x2; // @[MUL.scala 102:19]
  wire  m_1498_io_x3; // @[MUL.scala 102:19]
  wire  m_1498_io_s; // @[MUL.scala 102:19]
  wire  m_1498_io_cout; // @[MUL.scala 102:19]
  wire  m_1499_io_x1; // @[MUL.scala 102:19]
  wire  m_1499_io_x2; // @[MUL.scala 102:19]
  wire  m_1499_io_x3; // @[MUL.scala 102:19]
  wire  m_1499_io_s; // @[MUL.scala 102:19]
  wire  m_1499_io_cout; // @[MUL.scala 102:19]
  wire  m_1500_io_x1; // @[MUL.scala 102:19]
  wire  m_1500_io_x2; // @[MUL.scala 102:19]
  wire  m_1500_io_x3; // @[MUL.scala 102:19]
  wire  m_1500_io_s; // @[MUL.scala 102:19]
  wire  m_1500_io_cout; // @[MUL.scala 102:19]
  wire  m_1501_io_x1; // @[MUL.scala 102:19]
  wire  m_1501_io_x2; // @[MUL.scala 102:19]
  wire  m_1501_io_x3; // @[MUL.scala 102:19]
  wire  m_1501_io_s; // @[MUL.scala 102:19]
  wire  m_1501_io_cout; // @[MUL.scala 102:19]
  wire  m_1502_io_x1; // @[MUL.scala 102:19]
  wire  m_1502_io_x2; // @[MUL.scala 102:19]
  wire  m_1502_io_x3; // @[MUL.scala 102:19]
  wire  m_1502_io_s; // @[MUL.scala 102:19]
  wire  m_1502_io_cout; // @[MUL.scala 102:19]
  wire  m_1503_io_x1; // @[MUL.scala 102:19]
  wire  m_1503_io_x2; // @[MUL.scala 102:19]
  wire  m_1503_io_x3; // @[MUL.scala 102:19]
  wire  m_1503_io_s; // @[MUL.scala 102:19]
  wire  m_1503_io_cout; // @[MUL.scala 102:19]
  wire  m_1504_io_x1; // @[MUL.scala 102:19]
  wire  m_1504_io_x2; // @[MUL.scala 102:19]
  wire  m_1504_io_x3; // @[MUL.scala 102:19]
  wire  m_1504_io_s; // @[MUL.scala 102:19]
  wire  m_1504_io_cout; // @[MUL.scala 102:19]
  wire  m_1505_io_x1; // @[MUL.scala 102:19]
  wire  m_1505_io_x2; // @[MUL.scala 102:19]
  wire  m_1505_io_x3; // @[MUL.scala 102:19]
  wire  m_1505_io_s; // @[MUL.scala 102:19]
  wire  m_1505_io_cout; // @[MUL.scala 102:19]
  wire  m_1506_io_x1; // @[MUL.scala 102:19]
  wire  m_1506_io_x2; // @[MUL.scala 102:19]
  wire  m_1506_io_x3; // @[MUL.scala 102:19]
  wire  m_1506_io_s; // @[MUL.scala 102:19]
  wire  m_1506_io_cout; // @[MUL.scala 102:19]
  wire  m_1507_io_x1; // @[MUL.scala 102:19]
  wire  m_1507_io_x2; // @[MUL.scala 102:19]
  wire  m_1507_io_x3; // @[MUL.scala 102:19]
  wire  m_1507_io_s; // @[MUL.scala 102:19]
  wire  m_1507_io_cout; // @[MUL.scala 102:19]
  wire  m_1508_io_x1; // @[MUL.scala 102:19]
  wire  m_1508_io_x2; // @[MUL.scala 102:19]
  wire  m_1508_io_x3; // @[MUL.scala 102:19]
  wire  m_1508_io_s; // @[MUL.scala 102:19]
  wire  m_1508_io_cout; // @[MUL.scala 102:19]
  wire  m_1509_io_x1; // @[MUL.scala 102:19]
  wire  m_1509_io_x2; // @[MUL.scala 102:19]
  wire  m_1509_io_x3; // @[MUL.scala 102:19]
  wire  m_1509_io_s; // @[MUL.scala 102:19]
  wire  m_1509_io_cout; // @[MUL.scala 102:19]
  wire  m_1510_io_x1; // @[MUL.scala 102:19]
  wire  m_1510_io_x2; // @[MUL.scala 102:19]
  wire  m_1510_io_x3; // @[MUL.scala 102:19]
  wire  m_1510_io_s; // @[MUL.scala 102:19]
  wire  m_1510_io_cout; // @[MUL.scala 102:19]
  wire  m_1511_io_x1; // @[MUL.scala 102:19]
  wire  m_1511_io_x2; // @[MUL.scala 102:19]
  wire  m_1511_io_x3; // @[MUL.scala 102:19]
  wire  m_1511_io_s; // @[MUL.scala 102:19]
  wire  m_1511_io_cout; // @[MUL.scala 102:19]
  wire  m_1512_io_x1; // @[MUL.scala 102:19]
  wire  m_1512_io_x2; // @[MUL.scala 102:19]
  wire  m_1512_io_x3; // @[MUL.scala 102:19]
  wire  m_1512_io_s; // @[MUL.scala 102:19]
  wire  m_1512_io_cout; // @[MUL.scala 102:19]
  wire  m_1513_io_x1; // @[MUL.scala 102:19]
  wire  m_1513_io_x2; // @[MUL.scala 102:19]
  wire  m_1513_io_x3; // @[MUL.scala 102:19]
  wire  m_1513_io_s; // @[MUL.scala 102:19]
  wire  m_1513_io_cout; // @[MUL.scala 102:19]
  wire  m_1514_io_x1; // @[MUL.scala 102:19]
  wire  m_1514_io_x2; // @[MUL.scala 102:19]
  wire  m_1514_io_x3; // @[MUL.scala 102:19]
  wire  m_1514_io_s; // @[MUL.scala 102:19]
  wire  m_1514_io_cout; // @[MUL.scala 102:19]
  wire  m_1515_io_x1; // @[MUL.scala 102:19]
  wire  m_1515_io_x2; // @[MUL.scala 102:19]
  wire  m_1515_io_x3; // @[MUL.scala 102:19]
  wire  m_1515_io_s; // @[MUL.scala 102:19]
  wire  m_1515_io_cout; // @[MUL.scala 102:19]
  wire  m_1516_io_x1; // @[MUL.scala 102:19]
  wire  m_1516_io_x2; // @[MUL.scala 102:19]
  wire  m_1516_io_x3; // @[MUL.scala 102:19]
  wire  m_1516_io_s; // @[MUL.scala 102:19]
  wire  m_1516_io_cout; // @[MUL.scala 102:19]
  wire  m_1517_io_x1; // @[MUL.scala 102:19]
  wire  m_1517_io_x2; // @[MUL.scala 102:19]
  wire  m_1517_io_x3; // @[MUL.scala 102:19]
  wire  m_1517_io_s; // @[MUL.scala 102:19]
  wire  m_1517_io_cout; // @[MUL.scala 102:19]
  wire  m_1518_io_x1; // @[MUL.scala 102:19]
  wire  m_1518_io_x2; // @[MUL.scala 102:19]
  wire  m_1518_io_x3; // @[MUL.scala 102:19]
  wire  m_1518_io_s; // @[MUL.scala 102:19]
  wire  m_1518_io_cout; // @[MUL.scala 102:19]
  wire  m_1519_io_x1; // @[MUL.scala 102:19]
  wire  m_1519_io_x2; // @[MUL.scala 102:19]
  wire  m_1519_io_x3; // @[MUL.scala 102:19]
  wire  m_1519_io_s; // @[MUL.scala 102:19]
  wire  m_1519_io_cout; // @[MUL.scala 102:19]
  wire  m_1520_io_x1; // @[MUL.scala 102:19]
  wire  m_1520_io_x2; // @[MUL.scala 102:19]
  wire  m_1520_io_x3; // @[MUL.scala 102:19]
  wire  m_1520_io_s; // @[MUL.scala 102:19]
  wire  m_1520_io_cout; // @[MUL.scala 102:19]
  wire  m_1521_io_x1; // @[MUL.scala 102:19]
  wire  m_1521_io_x2; // @[MUL.scala 102:19]
  wire  m_1521_io_x3; // @[MUL.scala 102:19]
  wire  m_1521_io_s; // @[MUL.scala 102:19]
  wire  m_1521_io_cout; // @[MUL.scala 102:19]
  wire  m_1522_io_x1; // @[MUL.scala 102:19]
  wire  m_1522_io_x2; // @[MUL.scala 102:19]
  wire  m_1522_io_x3; // @[MUL.scala 102:19]
  wire  m_1522_io_s; // @[MUL.scala 102:19]
  wire  m_1522_io_cout; // @[MUL.scala 102:19]
  wire  m_1523_io_x1; // @[MUL.scala 102:19]
  wire  m_1523_io_x2; // @[MUL.scala 102:19]
  wire  m_1523_io_x3; // @[MUL.scala 102:19]
  wire  m_1523_io_s; // @[MUL.scala 102:19]
  wire  m_1523_io_cout; // @[MUL.scala 102:19]
  wire  m_1524_io_x1; // @[MUL.scala 102:19]
  wire  m_1524_io_x2; // @[MUL.scala 102:19]
  wire  m_1524_io_x3; // @[MUL.scala 102:19]
  wire  m_1524_io_s; // @[MUL.scala 102:19]
  wire  m_1524_io_cout; // @[MUL.scala 102:19]
  wire  m_1525_io_x1; // @[MUL.scala 102:19]
  wire  m_1525_io_x2; // @[MUL.scala 102:19]
  wire  m_1525_io_x3; // @[MUL.scala 102:19]
  wire  m_1525_io_s; // @[MUL.scala 102:19]
  wire  m_1525_io_cout; // @[MUL.scala 102:19]
  wire  m_1526_io_x1; // @[MUL.scala 102:19]
  wire  m_1526_io_x2; // @[MUL.scala 102:19]
  wire  m_1526_io_x3; // @[MUL.scala 102:19]
  wire  m_1526_io_s; // @[MUL.scala 102:19]
  wire  m_1526_io_cout; // @[MUL.scala 102:19]
  wire  m_1527_io_x1; // @[MUL.scala 102:19]
  wire  m_1527_io_x2; // @[MUL.scala 102:19]
  wire  m_1527_io_x3; // @[MUL.scala 102:19]
  wire  m_1527_io_s; // @[MUL.scala 102:19]
  wire  m_1527_io_cout; // @[MUL.scala 102:19]
  wire  m_1528_io_x1; // @[MUL.scala 102:19]
  wire  m_1528_io_x2; // @[MUL.scala 102:19]
  wire  m_1528_io_x3; // @[MUL.scala 102:19]
  wire  m_1528_io_s; // @[MUL.scala 102:19]
  wire  m_1528_io_cout; // @[MUL.scala 102:19]
  wire  m_1529_io_x1; // @[MUL.scala 102:19]
  wire  m_1529_io_x2; // @[MUL.scala 102:19]
  wire  m_1529_io_x3; // @[MUL.scala 102:19]
  wire  m_1529_io_s; // @[MUL.scala 102:19]
  wire  m_1529_io_cout; // @[MUL.scala 102:19]
  wire  m_1530_io_x1; // @[MUL.scala 102:19]
  wire  m_1530_io_x2; // @[MUL.scala 102:19]
  wire  m_1530_io_x3; // @[MUL.scala 102:19]
  wire  m_1530_io_s; // @[MUL.scala 102:19]
  wire  m_1530_io_cout; // @[MUL.scala 102:19]
  wire  m_1531_io_x1; // @[MUL.scala 102:19]
  wire  m_1531_io_x2; // @[MUL.scala 102:19]
  wire  m_1531_io_x3; // @[MUL.scala 102:19]
  wire  m_1531_io_s; // @[MUL.scala 102:19]
  wire  m_1531_io_cout; // @[MUL.scala 102:19]
  wire  m_1532_io_x1; // @[MUL.scala 102:19]
  wire  m_1532_io_x2; // @[MUL.scala 102:19]
  wire  m_1532_io_x3; // @[MUL.scala 102:19]
  wire  m_1532_io_s; // @[MUL.scala 102:19]
  wire  m_1532_io_cout; // @[MUL.scala 102:19]
  wire  m_1533_io_x1; // @[MUL.scala 102:19]
  wire  m_1533_io_x2; // @[MUL.scala 102:19]
  wire  m_1533_io_x3; // @[MUL.scala 102:19]
  wire  m_1533_io_s; // @[MUL.scala 102:19]
  wire  m_1533_io_cout; // @[MUL.scala 102:19]
  wire  m_1534_io_x1; // @[MUL.scala 102:19]
  wire  m_1534_io_x2; // @[MUL.scala 102:19]
  wire  m_1534_io_x3; // @[MUL.scala 102:19]
  wire  m_1534_io_s; // @[MUL.scala 102:19]
  wire  m_1534_io_cout; // @[MUL.scala 102:19]
  wire  m_1535_io_x1; // @[MUL.scala 102:19]
  wire  m_1535_io_x2; // @[MUL.scala 102:19]
  wire  m_1535_io_x3; // @[MUL.scala 102:19]
  wire  m_1535_io_s; // @[MUL.scala 102:19]
  wire  m_1535_io_cout; // @[MUL.scala 102:19]
  wire  m_1536_io_x1; // @[MUL.scala 102:19]
  wire  m_1536_io_x2; // @[MUL.scala 102:19]
  wire  m_1536_io_x3; // @[MUL.scala 102:19]
  wire  m_1536_io_s; // @[MUL.scala 102:19]
  wire  m_1536_io_cout; // @[MUL.scala 102:19]
  wire  m_1537_io_x1; // @[MUL.scala 102:19]
  wire  m_1537_io_x2; // @[MUL.scala 102:19]
  wire  m_1537_io_x3; // @[MUL.scala 102:19]
  wire  m_1537_io_s; // @[MUL.scala 102:19]
  wire  m_1537_io_cout; // @[MUL.scala 102:19]
  wire  m_1538_io_x1; // @[MUL.scala 102:19]
  wire  m_1538_io_x2; // @[MUL.scala 102:19]
  wire  m_1538_io_x3; // @[MUL.scala 102:19]
  wire  m_1538_io_s; // @[MUL.scala 102:19]
  wire  m_1538_io_cout; // @[MUL.scala 102:19]
  wire  m_1539_io_x1; // @[MUL.scala 102:19]
  wire  m_1539_io_x2; // @[MUL.scala 102:19]
  wire  m_1539_io_x3; // @[MUL.scala 102:19]
  wire  m_1539_io_s; // @[MUL.scala 102:19]
  wire  m_1539_io_cout; // @[MUL.scala 102:19]
  wire  m_1540_io_x1; // @[MUL.scala 102:19]
  wire  m_1540_io_x2; // @[MUL.scala 102:19]
  wire  m_1540_io_x3; // @[MUL.scala 102:19]
  wire  m_1540_io_s; // @[MUL.scala 102:19]
  wire  m_1540_io_cout; // @[MUL.scala 102:19]
  wire  m_1541_io_x1; // @[MUL.scala 102:19]
  wire  m_1541_io_x2; // @[MUL.scala 102:19]
  wire  m_1541_io_x3; // @[MUL.scala 102:19]
  wire  m_1541_io_s; // @[MUL.scala 102:19]
  wire  m_1541_io_cout; // @[MUL.scala 102:19]
  wire  m_1542_io_in_0; // @[MUL.scala 124:19]
  wire  m_1542_io_in_1; // @[MUL.scala 124:19]
  wire  m_1542_io_out_0; // @[MUL.scala 124:19]
  wire  m_1542_io_out_1; // @[MUL.scala 124:19]
  wire  m_1543_io_x1; // @[MUL.scala 102:19]
  wire  m_1543_io_x2; // @[MUL.scala 102:19]
  wire  m_1543_io_x3; // @[MUL.scala 102:19]
  wire  m_1543_io_s; // @[MUL.scala 102:19]
  wire  m_1543_io_cout; // @[MUL.scala 102:19]
  wire  m_1544_io_x1; // @[MUL.scala 102:19]
  wire  m_1544_io_x2; // @[MUL.scala 102:19]
  wire  m_1544_io_x3; // @[MUL.scala 102:19]
  wire  m_1544_io_s; // @[MUL.scala 102:19]
  wire  m_1544_io_cout; // @[MUL.scala 102:19]
  wire  m_1545_io_x1; // @[MUL.scala 102:19]
  wire  m_1545_io_x2; // @[MUL.scala 102:19]
  wire  m_1545_io_x3; // @[MUL.scala 102:19]
  wire  m_1545_io_s; // @[MUL.scala 102:19]
  wire  m_1545_io_cout; // @[MUL.scala 102:19]
  wire  m_1546_io_x1; // @[MUL.scala 102:19]
  wire  m_1546_io_x2; // @[MUL.scala 102:19]
  wire  m_1546_io_x3; // @[MUL.scala 102:19]
  wire  m_1546_io_s; // @[MUL.scala 102:19]
  wire  m_1546_io_cout; // @[MUL.scala 102:19]
  wire  m_1547_io_in_0; // @[MUL.scala 124:19]
  wire  m_1547_io_in_1; // @[MUL.scala 124:19]
  wire  m_1547_io_out_0; // @[MUL.scala 124:19]
  wire  m_1547_io_out_1; // @[MUL.scala 124:19]
  wire  m_1548_io_x1; // @[MUL.scala 102:19]
  wire  m_1548_io_x2; // @[MUL.scala 102:19]
  wire  m_1548_io_x3; // @[MUL.scala 102:19]
  wire  m_1548_io_s; // @[MUL.scala 102:19]
  wire  m_1548_io_cout; // @[MUL.scala 102:19]
  wire  m_1549_io_x1; // @[MUL.scala 102:19]
  wire  m_1549_io_x2; // @[MUL.scala 102:19]
  wire  m_1549_io_x3; // @[MUL.scala 102:19]
  wire  m_1549_io_s; // @[MUL.scala 102:19]
  wire  m_1549_io_cout; // @[MUL.scala 102:19]
  wire  m_1550_io_x1; // @[MUL.scala 102:19]
  wire  m_1550_io_x2; // @[MUL.scala 102:19]
  wire  m_1550_io_x3; // @[MUL.scala 102:19]
  wire  m_1550_io_s; // @[MUL.scala 102:19]
  wire  m_1550_io_cout; // @[MUL.scala 102:19]
  wire  m_1551_io_x1; // @[MUL.scala 102:19]
  wire  m_1551_io_x2; // @[MUL.scala 102:19]
  wire  m_1551_io_x3; // @[MUL.scala 102:19]
  wire  m_1551_io_s; // @[MUL.scala 102:19]
  wire  m_1551_io_cout; // @[MUL.scala 102:19]
  wire  m_1552_io_in_0; // @[MUL.scala 124:19]
  wire  m_1552_io_in_1; // @[MUL.scala 124:19]
  wire  m_1552_io_out_0; // @[MUL.scala 124:19]
  wire  m_1552_io_out_1; // @[MUL.scala 124:19]
  wire  m_1553_io_x1; // @[MUL.scala 102:19]
  wire  m_1553_io_x2; // @[MUL.scala 102:19]
  wire  m_1553_io_x3; // @[MUL.scala 102:19]
  wire  m_1553_io_s; // @[MUL.scala 102:19]
  wire  m_1553_io_cout; // @[MUL.scala 102:19]
  wire  m_1554_io_x1; // @[MUL.scala 102:19]
  wire  m_1554_io_x2; // @[MUL.scala 102:19]
  wire  m_1554_io_x3; // @[MUL.scala 102:19]
  wire  m_1554_io_s; // @[MUL.scala 102:19]
  wire  m_1554_io_cout; // @[MUL.scala 102:19]
  wire  m_1555_io_x1; // @[MUL.scala 102:19]
  wire  m_1555_io_x2; // @[MUL.scala 102:19]
  wire  m_1555_io_x3; // @[MUL.scala 102:19]
  wire  m_1555_io_s; // @[MUL.scala 102:19]
  wire  m_1555_io_cout; // @[MUL.scala 102:19]
  wire  m_1556_io_x1; // @[MUL.scala 102:19]
  wire  m_1556_io_x2; // @[MUL.scala 102:19]
  wire  m_1556_io_x3; // @[MUL.scala 102:19]
  wire  m_1556_io_s; // @[MUL.scala 102:19]
  wire  m_1556_io_cout; // @[MUL.scala 102:19]
  wire  m_1557_io_in_0; // @[MUL.scala 124:19]
  wire  m_1557_io_in_1; // @[MUL.scala 124:19]
  wire  m_1557_io_out_0; // @[MUL.scala 124:19]
  wire  m_1557_io_out_1; // @[MUL.scala 124:19]
  wire  m_1558_io_x1; // @[MUL.scala 102:19]
  wire  m_1558_io_x2; // @[MUL.scala 102:19]
  wire  m_1558_io_x3; // @[MUL.scala 102:19]
  wire  m_1558_io_s; // @[MUL.scala 102:19]
  wire  m_1558_io_cout; // @[MUL.scala 102:19]
  wire  m_1559_io_x1; // @[MUL.scala 102:19]
  wire  m_1559_io_x2; // @[MUL.scala 102:19]
  wire  m_1559_io_x3; // @[MUL.scala 102:19]
  wire  m_1559_io_s; // @[MUL.scala 102:19]
  wire  m_1559_io_cout; // @[MUL.scala 102:19]
  wire  m_1560_io_x1; // @[MUL.scala 102:19]
  wire  m_1560_io_x2; // @[MUL.scala 102:19]
  wire  m_1560_io_x3; // @[MUL.scala 102:19]
  wire  m_1560_io_s; // @[MUL.scala 102:19]
  wire  m_1560_io_cout; // @[MUL.scala 102:19]
  wire  m_1561_io_x1; // @[MUL.scala 102:19]
  wire  m_1561_io_x2; // @[MUL.scala 102:19]
  wire  m_1561_io_x3; // @[MUL.scala 102:19]
  wire  m_1561_io_s; // @[MUL.scala 102:19]
  wire  m_1561_io_cout; // @[MUL.scala 102:19]
  wire  m_1562_io_in_0; // @[MUL.scala 124:19]
  wire  m_1562_io_in_1; // @[MUL.scala 124:19]
  wire  m_1562_io_out_0; // @[MUL.scala 124:19]
  wire  m_1562_io_out_1; // @[MUL.scala 124:19]
  wire  m_1563_io_x1; // @[MUL.scala 102:19]
  wire  m_1563_io_x2; // @[MUL.scala 102:19]
  wire  m_1563_io_x3; // @[MUL.scala 102:19]
  wire  m_1563_io_s; // @[MUL.scala 102:19]
  wire  m_1563_io_cout; // @[MUL.scala 102:19]
  wire  m_1564_io_x1; // @[MUL.scala 102:19]
  wire  m_1564_io_x2; // @[MUL.scala 102:19]
  wire  m_1564_io_x3; // @[MUL.scala 102:19]
  wire  m_1564_io_s; // @[MUL.scala 102:19]
  wire  m_1564_io_cout; // @[MUL.scala 102:19]
  wire  m_1565_io_x1; // @[MUL.scala 102:19]
  wire  m_1565_io_x2; // @[MUL.scala 102:19]
  wire  m_1565_io_x3; // @[MUL.scala 102:19]
  wire  m_1565_io_s; // @[MUL.scala 102:19]
  wire  m_1565_io_cout; // @[MUL.scala 102:19]
  wire  m_1566_io_x1; // @[MUL.scala 102:19]
  wire  m_1566_io_x2; // @[MUL.scala 102:19]
  wire  m_1566_io_x3; // @[MUL.scala 102:19]
  wire  m_1566_io_s; // @[MUL.scala 102:19]
  wire  m_1566_io_cout; // @[MUL.scala 102:19]
  wire  m_1567_io_in_0; // @[MUL.scala 124:19]
  wire  m_1567_io_in_1; // @[MUL.scala 124:19]
  wire  m_1567_io_out_0; // @[MUL.scala 124:19]
  wire  m_1567_io_out_1; // @[MUL.scala 124:19]
  wire  m_1568_io_x1; // @[MUL.scala 102:19]
  wire  m_1568_io_x2; // @[MUL.scala 102:19]
  wire  m_1568_io_x3; // @[MUL.scala 102:19]
  wire  m_1568_io_s; // @[MUL.scala 102:19]
  wire  m_1568_io_cout; // @[MUL.scala 102:19]
  wire  m_1569_io_x1; // @[MUL.scala 102:19]
  wire  m_1569_io_x2; // @[MUL.scala 102:19]
  wire  m_1569_io_x3; // @[MUL.scala 102:19]
  wire  m_1569_io_s; // @[MUL.scala 102:19]
  wire  m_1569_io_cout; // @[MUL.scala 102:19]
  wire  m_1570_io_x1; // @[MUL.scala 102:19]
  wire  m_1570_io_x2; // @[MUL.scala 102:19]
  wire  m_1570_io_x3; // @[MUL.scala 102:19]
  wire  m_1570_io_s; // @[MUL.scala 102:19]
  wire  m_1570_io_cout; // @[MUL.scala 102:19]
  wire  m_1571_io_x1; // @[MUL.scala 102:19]
  wire  m_1571_io_x2; // @[MUL.scala 102:19]
  wire  m_1571_io_x3; // @[MUL.scala 102:19]
  wire  m_1571_io_s; // @[MUL.scala 102:19]
  wire  m_1571_io_cout; // @[MUL.scala 102:19]
  wire  m_1572_io_in_0; // @[MUL.scala 124:19]
  wire  m_1572_io_in_1; // @[MUL.scala 124:19]
  wire  m_1572_io_out_0; // @[MUL.scala 124:19]
  wire  m_1572_io_out_1; // @[MUL.scala 124:19]
  wire  m_1573_io_x1; // @[MUL.scala 102:19]
  wire  m_1573_io_x2; // @[MUL.scala 102:19]
  wire  m_1573_io_x3; // @[MUL.scala 102:19]
  wire  m_1573_io_s; // @[MUL.scala 102:19]
  wire  m_1573_io_cout; // @[MUL.scala 102:19]
  wire  m_1574_io_x1; // @[MUL.scala 102:19]
  wire  m_1574_io_x2; // @[MUL.scala 102:19]
  wire  m_1574_io_x3; // @[MUL.scala 102:19]
  wire  m_1574_io_s; // @[MUL.scala 102:19]
  wire  m_1574_io_cout; // @[MUL.scala 102:19]
  wire  m_1575_io_x1; // @[MUL.scala 102:19]
  wire  m_1575_io_x2; // @[MUL.scala 102:19]
  wire  m_1575_io_x3; // @[MUL.scala 102:19]
  wire  m_1575_io_s; // @[MUL.scala 102:19]
  wire  m_1575_io_cout; // @[MUL.scala 102:19]
  wire  m_1576_io_x1; // @[MUL.scala 102:19]
  wire  m_1576_io_x2; // @[MUL.scala 102:19]
  wire  m_1576_io_x3; // @[MUL.scala 102:19]
  wire  m_1576_io_s; // @[MUL.scala 102:19]
  wire  m_1576_io_cout; // @[MUL.scala 102:19]
  wire  m_1577_io_x1; // @[MUL.scala 102:19]
  wire  m_1577_io_x2; // @[MUL.scala 102:19]
  wire  m_1577_io_x3; // @[MUL.scala 102:19]
  wire  m_1577_io_s; // @[MUL.scala 102:19]
  wire  m_1577_io_cout; // @[MUL.scala 102:19]
  wire  m_1578_io_x1; // @[MUL.scala 102:19]
  wire  m_1578_io_x2; // @[MUL.scala 102:19]
  wire  m_1578_io_x3; // @[MUL.scala 102:19]
  wire  m_1578_io_s; // @[MUL.scala 102:19]
  wire  m_1578_io_cout; // @[MUL.scala 102:19]
  wire  m_1579_io_x1; // @[MUL.scala 102:19]
  wire  m_1579_io_x2; // @[MUL.scala 102:19]
  wire  m_1579_io_x3; // @[MUL.scala 102:19]
  wire  m_1579_io_s; // @[MUL.scala 102:19]
  wire  m_1579_io_cout; // @[MUL.scala 102:19]
  wire  m_1580_io_x1; // @[MUL.scala 102:19]
  wire  m_1580_io_x2; // @[MUL.scala 102:19]
  wire  m_1580_io_x3; // @[MUL.scala 102:19]
  wire  m_1580_io_s; // @[MUL.scala 102:19]
  wire  m_1580_io_cout; // @[MUL.scala 102:19]
  wire  m_1581_io_x1; // @[MUL.scala 102:19]
  wire  m_1581_io_x2; // @[MUL.scala 102:19]
  wire  m_1581_io_x3; // @[MUL.scala 102:19]
  wire  m_1581_io_s; // @[MUL.scala 102:19]
  wire  m_1581_io_cout; // @[MUL.scala 102:19]
  wire  m_1582_io_x1; // @[MUL.scala 102:19]
  wire  m_1582_io_x2; // @[MUL.scala 102:19]
  wire  m_1582_io_x3; // @[MUL.scala 102:19]
  wire  m_1582_io_s; // @[MUL.scala 102:19]
  wire  m_1582_io_cout; // @[MUL.scala 102:19]
  wire  m_1583_io_x1; // @[MUL.scala 102:19]
  wire  m_1583_io_x2; // @[MUL.scala 102:19]
  wire  m_1583_io_x3; // @[MUL.scala 102:19]
  wire  m_1583_io_s; // @[MUL.scala 102:19]
  wire  m_1583_io_cout; // @[MUL.scala 102:19]
  wire  m_1584_io_x1; // @[MUL.scala 102:19]
  wire  m_1584_io_x2; // @[MUL.scala 102:19]
  wire  m_1584_io_x3; // @[MUL.scala 102:19]
  wire  m_1584_io_s; // @[MUL.scala 102:19]
  wire  m_1584_io_cout; // @[MUL.scala 102:19]
  wire  m_1585_io_x1; // @[MUL.scala 102:19]
  wire  m_1585_io_x2; // @[MUL.scala 102:19]
  wire  m_1585_io_x3; // @[MUL.scala 102:19]
  wire  m_1585_io_s; // @[MUL.scala 102:19]
  wire  m_1585_io_cout; // @[MUL.scala 102:19]
  wire  m_1586_io_x1; // @[MUL.scala 102:19]
  wire  m_1586_io_x2; // @[MUL.scala 102:19]
  wire  m_1586_io_x3; // @[MUL.scala 102:19]
  wire  m_1586_io_s; // @[MUL.scala 102:19]
  wire  m_1586_io_cout; // @[MUL.scala 102:19]
  wire  m_1587_io_x1; // @[MUL.scala 102:19]
  wire  m_1587_io_x2; // @[MUL.scala 102:19]
  wire  m_1587_io_x3; // @[MUL.scala 102:19]
  wire  m_1587_io_s; // @[MUL.scala 102:19]
  wire  m_1587_io_cout; // @[MUL.scala 102:19]
  wire  m_1588_io_x1; // @[MUL.scala 102:19]
  wire  m_1588_io_x2; // @[MUL.scala 102:19]
  wire  m_1588_io_x3; // @[MUL.scala 102:19]
  wire  m_1588_io_s; // @[MUL.scala 102:19]
  wire  m_1588_io_cout; // @[MUL.scala 102:19]
  wire  m_1589_io_x1; // @[MUL.scala 102:19]
  wire  m_1589_io_x2; // @[MUL.scala 102:19]
  wire  m_1589_io_x3; // @[MUL.scala 102:19]
  wire  m_1589_io_s; // @[MUL.scala 102:19]
  wire  m_1589_io_cout; // @[MUL.scala 102:19]
  wire  m_1590_io_x1; // @[MUL.scala 102:19]
  wire  m_1590_io_x2; // @[MUL.scala 102:19]
  wire  m_1590_io_x3; // @[MUL.scala 102:19]
  wire  m_1590_io_s; // @[MUL.scala 102:19]
  wire  m_1590_io_cout; // @[MUL.scala 102:19]
  wire  m_1591_io_x1; // @[MUL.scala 102:19]
  wire  m_1591_io_x2; // @[MUL.scala 102:19]
  wire  m_1591_io_x3; // @[MUL.scala 102:19]
  wire  m_1591_io_s; // @[MUL.scala 102:19]
  wire  m_1591_io_cout; // @[MUL.scala 102:19]
  wire  m_1592_io_x1; // @[MUL.scala 102:19]
  wire  m_1592_io_x2; // @[MUL.scala 102:19]
  wire  m_1592_io_x3; // @[MUL.scala 102:19]
  wire  m_1592_io_s; // @[MUL.scala 102:19]
  wire  m_1592_io_cout; // @[MUL.scala 102:19]
  wire  m_1593_io_x1; // @[MUL.scala 102:19]
  wire  m_1593_io_x2; // @[MUL.scala 102:19]
  wire  m_1593_io_x3; // @[MUL.scala 102:19]
  wire  m_1593_io_s; // @[MUL.scala 102:19]
  wire  m_1593_io_cout; // @[MUL.scala 102:19]
  wire  m_1594_io_x1; // @[MUL.scala 102:19]
  wire  m_1594_io_x2; // @[MUL.scala 102:19]
  wire  m_1594_io_x3; // @[MUL.scala 102:19]
  wire  m_1594_io_s; // @[MUL.scala 102:19]
  wire  m_1594_io_cout; // @[MUL.scala 102:19]
  wire  m_1595_io_x1; // @[MUL.scala 102:19]
  wire  m_1595_io_x2; // @[MUL.scala 102:19]
  wire  m_1595_io_x3; // @[MUL.scala 102:19]
  wire  m_1595_io_s; // @[MUL.scala 102:19]
  wire  m_1595_io_cout; // @[MUL.scala 102:19]
  wire  m_1596_io_x1; // @[MUL.scala 102:19]
  wire  m_1596_io_x2; // @[MUL.scala 102:19]
  wire  m_1596_io_x3; // @[MUL.scala 102:19]
  wire  m_1596_io_s; // @[MUL.scala 102:19]
  wire  m_1596_io_cout; // @[MUL.scala 102:19]
  wire  m_1597_io_x1; // @[MUL.scala 102:19]
  wire  m_1597_io_x2; // @[MUL.scala 102:19]
  wire  m_1597_io_x3; // @[MUL.scala 102:19]
  wire  m_1597_io_s; // @[MUL.scala 102:19]
  wire  m_1597_io_cout; // @[MUL.scala 102:19]
  wire  m_1598_io_x1; // @[MUL.scala 102:19]
  wire  m_1598_io_x2; // @[MUL.scala 102:19]
  wire  m_1598_io_x3; // @[MUL.scala 102:19]
  wire  m_1598_io_s; // @[MUL.scala 102:19]
  wire  m_1598_io_cout; // @[MUL.scala 102:19]
  wire  m_1599_io_x1; // @[MUL.scala 102:19]
  wire  m_1599_io_x2; // @[MUL.scala 102:19]
  wire  m_1599_io_x3; // @[MUL.scala 102:19]
  wire  m_1599_io_s; // @[MUL.scala 102:19]
  wire  m_1599_io_cout; // @[MUL.scala 102:19]
  wire  m_1600_io_x1; // @[MUL.scala 102:19]
  wire  m_1600_io_x2; // @[MUL.scala 102:19]
  wire  m_1600_io_x3; // @[MUL.scala 102:19]
  wire  m_1600_io_s; // @[MUL.scala 102:19]
  wire  m_1600_io_cout; // @[MUL.scala 102:19]
  wire  m_1601_io_x1; // @[MUL.scala 102:19]
  wire  m_1601_io_x2; // @[MUL.scala 102:19]
  wire  m_1601_io_x3; // @[MUL.scala 102:19]
  wire  m_1601_io_s; // @[MUL.scala 102:19]
  wire  m_1601_io_cout; // @[MUL.scala 102:19]
  wire  m_1602_io_x1; // @[MUL.scala 102:19]
  wire  m_1602_io_x2; // @[MUL.scala 102:19]
  wire  m_1602_io_x3; // @[MUL.scala 102:19]
  wire  m_1602_io_s; // @[MUL.scala 102:19]
  wire  m_1602_io_cout; // @[MUL.scala 102:19]
  wire  m_1603_io_x1; // @[MUL.scala 102:19]
  wire  m_1603_io_x2; // @[MUL.scala 102:19]
  wire  m_1603_io_x3; // @[MUL.scala 102:19]
  wire  m_1603_io_s; // @[MUL.scala 102:19]
  wire  m_1603_io_cout; // @[MUL.scala 102:19]
  wire  m_1604_io_in_0; // @[MUL.scala 124:19]
  wire  m_1604_io_in_1; // @[MUL.scala 124:19]
  wire  m_1604_io_out_0; // @[MUL.scala 124:19]
  wire  m_1604_io_out_1; // @[MUL.scala 124:19]
  wire  m_1605_io_x1; // @[MUL.scala 102:19]
  wire  m_1605_io_x2; // @[MUL.scala 102:19]
  wire  m_1605_io_x3; // @[MUL.scala 102:19]
  wire  m_1605_io_s; // @[MUL.scala 102:19]
  wire  m_1605_io_cout; // @[MUL.scala 102:19]
  wire  m_1606_io_x1; // @[MUL.scala 102:19]
  wire  m_1606_io_x2; // @[MUL.scala 102:19]
  wire  m_1606_io_x3; // @[MUL.scala 102:19]
  wire  m_1606_io_s; // @[MUL.scala 102:19]
  wire  m_1606_io_cout; // @[MUL.scala 102:19]
  wire  m_1607_io_x1; // @[MUL.scala 102:19]
  wire  m_1607_io_x2; // @[MUL.scala 102:19]
  wire  m_1607_io_x3; // @[MUL.scala 102:19]
  wire  m_1607_io_s; // @[MUL.scala 102:19]
  wire  m_1607_io_cout; // @[MUL.scala 102:19]
  wire  m_1608_io_in_0; // @[MUL.scala 124:19]
  wire  m_1608_io_in_1; // @[MUL.scala 124:19]
  wire  m_1608_io_out_0; // @[MUL.scala 124:19]
  wire  m_1608_io_out_1; // @[MUL.scala 124:19]
  wire  m_1609_io_x1; // @[MUL.scala 102:19]
  wire  m_1609_io_x2; // @[MUL.scala 102:19]
  wire  m_1609_io_x3; // @[MUL.scala 102:19]
  wire  m_1609_io_s; // @[MUL.scala 102:19]
  wire  m_1609_io_cout; // @[MUL.scala 102:19]
  wire  m_1610_io_x1; // @[MUL.scala 102:19]
  wire  m_1610_io_x2; // @[MUL.scala 102:19]
  wire  m_1610_io_x3; // @[MUL.scala 102:19]
  wire  m_1610_io_s; // @[MUL.scala 102:19]
  wire  m_1610_io_cout; // @[MUL.scala 102:19]
  wire  m_1611_io_x1; // @[MUL.scala 102:19]
  wire  m_1611_io_x2; // @[MUL.scala 102:19]
  wire  m_1611_io_x3; // @[MUL.scala 102:19]
  wire  m_1611_io_s; // @[MUL.scala 102:19]
  wire  m_1611_io_cout; // @[MUL.scala 102:19]
  wire  m_1612_io_in_0; // @[MUL.scala 124:19]
  wire  m_1612_io_in_1; // @[MUL.scala 124:19]
  wire  m_1612_io_out_0; // @[MUL.scala 124:19]
  wire  m_1612_io_out_1; // @[MUL.scala 124:19]
  wire  m_1613_io_x1; // @[MUL.scala 102:19]
  wire  m_1613_io_x2; // @[MUL.scala 102:19]
  wire  m_1613_io_x3; // @[MUL.scala 102:19]
  wire  m_1613_io_s; // @[MUL.scala 102:19]
  wire  m_1613_io_cout; // @[MUL.scala 102:19]
  wire  m_1614_io_x1; // @[MUL.scala 102:19]
  wire  m_1614_io_x2; // @[MUL.scala 102:19]
  wire  m_1614_io_x3; // @[MUL.scala 102:19]
  wire  m_1614_io_s; // @[MUL.scala 102:19]
  wire  m_1614_io_cout; // @[MUL.scala 102:19]
  wire  m_1615_io_x1; // @[MUL.scala 102:19]
  wire  m_1615_io_x2; // @[MUL.scala 102:19]
  wire  m_1615_io_x3; // @[MUL.scala 102:19]
  wire  m_1615_io_s; // @[MUL.scala 102:19]
  wire  m_1615_io_cout; // @[MUL.scala 102:19]
  wire  m_1616_io_in_0; // @[MUL.scala 124:19]
  wire  m_1616_io_in_1; // @[MUL.scala 124:19]
  wire  m_1616_io_out_0; // @[MUL.scala 124:19]
  wire  m_1616_io_out_1; // @[MUL.scala 124:19]
  wire  m_1617_io_x1; // @[MUL.scala 102:19]
  wire  m_1617_io_x2; // @[MUL.scala 102:19]
  wire  m_1617_io_x3; // @[MUL.scala 102:19]
  wire  m_1617_io_s; // @[MUL.scala 102:19]
  wire  m_1617_io_cout; // @[MUL.scala 102:19]
  wire  m_1618_io_x1; // @[MUL.scala 102:19]
  wire  m_1618_io_x2; // @[MUL.scala 102:19]
  wire  m_1618_io_x3; // @[MUL.scala 102:19]
  wire  m_1618_io_s; // @[MUL.scala 102:19]
  wire  m_1618_io_cout; // @[MUL.scala 102:19]
  wire  m_1619_io_x1; // @[MUL.scala 102:19]
  wire  m_1619_io_x2; // @[MUL.scala 102:19]
  wire  m_1619_io_x3; // @[MUL.scala 102:19]
  wire  m_1619_io_s; // @[MUL.scala 102:19]
  wire  m_1619_io_cout; // @[MUL.scala 102:19]
  wire  m_1620_io_x1; // @[MUL.scala 102:19]
  wire  m_1620_io_x2; // @[MUL.scala 102:19]
  wire  m_1620_io_x3; // @[MUL.scala 102:19]
  wire  m_1620_io_s; // @[MUL.scala 102:19]
  wire  m_1620_io_cout; // @[MUL.scala 102:19]
  wire  m_1621_io_x1; // @[MUL.scala 102:19]
  wire  m_1621_io_x2; // @[MUL.scala 102:19]
  wire  m_1621_io_x3; // @[MUL.scala 102:19]
  wire  m_1621_io_s; // @[MUL.scala 102:19]
  wire  m_1621_io_cout; // @[MUL.scala 102:19]
  wire  m_1622_io_x1; // @[MUL.scala 102:19]
  wire  m_1622_io_x2; // @[MUL.scala 102:19]
  wire  m_1622_io_x3; // @[MUL.scala 102:19]
  wire  m_1622_io_s; // @[MUL.scala 102:19]
  wire  m_1622_io_cout; // @[MUL.scala 102:19]
  wire  m_1623_io_x1; // @[MUL.scala 102:19]
  wire  m_1623_io_x2; // @[MUL.scala 102:19]
  wire  m_1623_io_x3; // @[MUL.scala 102:19]
  wire  m_1623_io_s; // @[MUL.scala 102:19]
  wire  m_1623_io_cout; // @[MUL.scala 102:19]
  wire  m_1624_io_x1; // @[MUL.scala 102:19]
  wire  m_1624_io_x2; // @[MUL.scala 102:19]
  wire  m_1624_io_x3; // @[MUL.scala 102:19]
  wire  m_1624_io_s; // @[MUL.scala 102:19]
  wire  m_1624_io_cout; // @[MUL.scala 102:19]
  wire  m_1625_io_x1; // @[MUL.scala 102:19]
  wire  m_1625_io_x2; // @[MUL.scala 102:19]
  wire  m_1625_io_x3; // @[MUL.scala 102:19]
  wire  m_1625_io_s; // @[MUL.scala 102:19]
  wire  m_1625_io_cout; // @[MUL.scala 102:19]
  wire  m_1626_io_x1; // @[MUL.scala 102:19]
  wire  m_1626_io_x2; // @[MUL.scala 102:19]
  wire  m_1626_io_x3; // @[MUL.scala 102:19]
  wire  m_1626_io_s; // @[MUL.scala 102:19]
  wire  m_1626_io_cout; // @[MUL.scala 102:19]
  wire  m_1627_io_x1; // @[MUL.scala 102:19]
  wire  m_1627_io_x2; // @[MUL.scala 102:19]
  wire  m_1627_io_x3; // @[MUL.scala 102:19]
  wire  m_1627_io_s; // @[MUL.scala 102:19]
  wire  m_1627_io_cout; // @[MUL.scala 102:19]
  wire  m_1628_io_x1; // @[MUL.scala 102:19]
  wire  m_1628_io_x2; // @[MUL.scala 102:19]
  wire  m_1628_io_x3; // @[MUL.scala 102:19]
  wire  m_1628_io_s; // @[MUL.scala 102:19]
  wire  m_1628_io_cout; // @[MUL.scala 102:19]
  wire  m_1629_io_x1; // @[MUL.scala 102:19]
  wire  m_1629_io_x2; // @[MUL.scala 102:19]
  wire  m_1629_io_x3; // @[MUL.scala 102:19]
  wire  m_1629_io_s; // @[MUL.scala 102:19]
  wire  m_1629_io_cout; // @[MUL.scala 102:19]
  wire  m_1630_io_x1; // @[MUL.scala 102:19]
  wire  m_1630_io_x2; // @[MUL.scala 102:19]
  wire  m_1630_io_x3; // @[MUL.scala 102:19]
  wire  m_1630_io_s; // @[MUL.scala 102:19]
  wire  m_1630_io_cout; // @[MUL.scala 102:19]
  wire  m_1631_io_x1; // @[MUL.scala 102:19]
  wire  m_1631_io_x2; // @[MUL.scala 102:19]
  wire  m_1631_io_x3; // @[MUL.scala 102:19]
  wire  m_1631_io_s; // @[MUL.scala 102:19]
  wire  m_1631_io_cout; // @[MUL.scala 102:19]
  wire  m_1632_io_x1; // @[MUL.scala 102:19]
  wire  m_1632_io_x2; // @[MUL.scala 102:19]
  wire  m_1632_io_x3; // @[MUL.scala 102:19]
  wire  m_1632_io_s; // @[MUL.scala 102:19]
  wire  m_1632_io_cout; // @[MUL.scala 102:19]
  wire  m_1633_io_x1; // @[MUL.scala 102:19]
  wire  m_1633_io_x2; // @[MUL.scala 102:19]
  wire  m_1633_io_x3; // @[MUL.scala 102:19]
  wire  m_1633_io_s; // @[MUL.scala 102:19]
  wire  m_1633_io_cout; // @[MUL.scala 102:19]
  wire  m_1634_io_x1; // @[MUL.scala 102:19]
  wire  m_1634_io_x2; // @[MUL.scala 102:19]
  wire  m_1634_io_x3; // @[MUL.scala 102:19]
  wire  m_1634_io_s; // @[MUL.scala 102:19]
  wire  m_1634_io_cout; // @[MUL.scala 102:19]
  wire  m_1635_io_x1; // @[MUL.scala 102:19]
  wire  m_1635_io_x2; // @[MUL.scala 102:19]
  wire  m_1635_io_x3; // @[MUL.scala 102:19]
  wire  m_1635_io_s; // @[MUL.scala 102:19]
  wire  m_1635_io_cout; // @[MUL.scala 102:19]
  wire  m_1636_io_x1; // @[MUL.scala 102:19]
  wire  m_1636_io_x2; // @[MUL.scala 102:19]
  wire  m_1636_io_x3; // @[MUL.scala 102:19]
  wire  m_1636_io_s; // @[MUL.scala 102:19]
  wire  m_1636_io_cout; // @[MUL.scala 102:19]
  wire  m_1637_io_x1; // @[MUL.scala 102:19]
  wire  m_1637_io_x2; // @[MUL.scala 102:19]
  wire  m_1637_io_x3; // @[MUL.scala 102:19]
  wire  m_1637_io_s; // @[MUL.scala 102:19]
  wire  m_1637_io_cout; // @[MUL.scala 102:19]
  wire  m_1638_io_x1; // @[MUL.scala 102:19]
  wire  m_1638_io_x2; // @[MUL.scala 102:19]
  wire  m_1638_io_x3; // @[MUL.scala 102:19]
  wire  m_1638_io_s; // @[MUL.scala 102:19]
  wire  m_1638_io_cout; // @[MUL.scala 102:19]
  wire  m_1639_io_x1; // @[MUL.scala 102:19]
  wire  m_1639_io_x2; // @[MUL.scala 102:19]
  wire  m_1639_io_x3; // @[MUL.scala 102:19]
  wire  m_1639_io_s; // @[MUL.scala 102:19]
  wire  m_1639_io_cout; // @[MUL.scala 102:19]
  wire  m_1640_io_in_0; // @[MUL.scala 124:19]
  wire  m_1640_io_in_1; // @[MUL.scala 124:19]
  wire  m_1640_io_out_0; // @[MUL.scala 124:19]
  wire  m_1640_io_out_1; // @[MUL.scala 124:19]
  wire  m_1641_io_x1; // @[MUL.scala 102:19]
  wire  m_1641_io_x2; // @[MUL.scala 102:19]
  wire  m_1641_io_x3; // @[MUL.scala 102:19]
  wire  m_1641_io_s; // @[MUL.scala 102:19]
  wire  m_1641_io_cout; // @[MUL.scala 102:19]
  wire  m_1642_io_x1; // @[MUL.scala 102:19]
  wire  m_1642_io_x2; // @[MUL.scala 102:19]
  wire  m_1642_io_x3; // @[MUL.scala 102:19]
  wire  m_1642_io_s; // @[MUL.scala 102:19]
  wire  m_1642_io_cout; // @[MUL.scala 102:19]
  wire  m_1643_io_in_0; // @[MUL.scala 124:19]
  wire  m_1643_io_in_1; // @[MUL.scala 124:19]
  wire  m_1643_io_out_0; // @[MUL.scala 124:19]
  wire  m_1643_io_out_1; // @[MUL.scala 124:19]
  wire  m_1644_io_x1; // @[MUL.scala 102:19]
  wire  m_1644_io_x2; // @[MUL.scala 102:19]
  wire  m_1644_io_x3; // @[MUL.scala 102:19]
  wire  m_1644_io_s; // @[MUL.scala 102:19]
  wire  m_1644_io_cout; // @[MUL.scala 102:19]
  wire  m_1645_io_x1; // @[MUL.scala 102:19]
  wire  m_1645_io_x2; // @[MUL.scala 102:19]
  wire  m_1645_io_x3; // @[MUL.scala 102:19]
  wire  m_1645_io_s; // @[MUL.scala 102:19]
  wire  m_1645_io_cout; // @[MUL.scala 102:19]
  wire  m_1646_io_in_0; // @[MUL.scala 124:19]
  wire  m_1646_io_in_1; // @[MUL.scala 124:19]
  wire  m_1646_io_out_0; // @[MUL.scala 124:19]
  wire  m_1646_io_out_1; // @[MUL.scala 124:19]
  wire  m_1647_io_x1; // @[MUL.scala 102:19]
  wire  m_1647_io_x2; // @[MUL.scala 102:19]
  wire  m_1647_io_x3; // @[MUL.scala 102:19]
  wire  m_1647_io_s; // @[MUL.scala 102:19]
  wire  m_1647_io_cout; // @[MUL.scala 102:19]
  wire  m_1648_io_x1; // @[MUL.scala 102:19]
  wire  m_1648_io_x2; // @[MUL.scala 102:19]
  wire  m_1648_io_x3; // @[MUL.scala 102:19]
  wire  m_1648_io_s; // @[MUL.scala 102:19]
  wire  m_1648_io_cout; // @[MUL.scala 102:19]
  wire  m_1649_io_in_0; // @[MUL.scala 124:19]
  wire  m_1649_io_in_1; // @[MUL.scala 124:19]
  wire  m_1649_io_out_0; // @[MUL.scala 124:19]
  wire  m_1649_io_out_1; // @[MUL.scala 124:19]
  wire  m_1650_io_x1; // @[MUL.scala 102:19]
  wire  m_1650_io_x2; // @[MUL.scala 102:19]
  wire  m_1650_io_x3; // @[MUL.scala 102:19]
  wire  m_1650_io_s; // @[MUL.scala 102:19]
  wire  m_1650_io_cout; // @[MUL.scala 102:19]
  wire  m_1651_io_x1; // @[MUL.scala 102:19]
  wire  m_1651_io_x2; // @[MUL.scala 102:19]
  wire  m_1651_io_x3; // @[MUL.scala 102:19]
  wire  m_1651_io_s; // @[MUL.scala 102:19]
  wire  m_1651_io_cout; // @[MUL.scala 102:19]
  wire  m_1652_io_in_0; // @[MUL.scala 124:19]
  wire  m_1652_io_in_1; // @[MUL.scala 124:19]
  wire  m_1652_io_out_0; // @[MUL.scala 124:19]
  wire  m_1652_io_out_1; // @[MUL.scala 124:19]
  wire  m_1653_io_x1; // @[MUL.scala 102:19]
  wire  m_1653_io_x2; // @[MUL.scala 102:19]
  wire  m_1653_io_x3; // @[MUL.scala 102:19]
  wire  m_1653_io_s; // @[MUL.scala 102:19]
  wire  m_1653_io_cout; // @[MUL.scala 102:19]
  wire  m_1654_io_x1; // @[MUL.scala 102:19]
  wire  m_1654_io_x2; // @[MUL.scala 102:19]
  wire  m_1654_io_x3; // @[MUL.scala 102:19]
  wire  m_1654_io_s; // @[MUL.scala 102:19]
  wire  m_1654_io_cout; // @[MUL.scala 102:19]
  wire  m_1655_io_in_0; // @[MUL.scala 124:19]
  wire  m_1655_io_in_1; // @[MUL.scala 124:19]
  wire  m_1655_io_out_0; // @[MUL.scala 124:19]
  wire  m_1655_io_out_1; // @[MUL.scala 124:19]
  wire  m_1656_io_x1; // @[MUL.scala 102:19]
  wire  m_1656_io_x2; // @[MUL.scala 102:19]
  wire  m_1656_io_x3; // @[MUL.scala 102:19]
  wire  m_1656_io_s; // @[MUL.scala 102:19]
  wire  m_1656_io_cout; // @[MUL.scala 102:19]
  wire  m_1657_io_x1; // @[MUL.scala 102:19]
  wire  m_1657_io_x2; // @[MUL.scala 102:19]
  wire  m_1657_io_x3; // @[MUL.scala 102:19]
  wire  m_1657_io_s; // @[MUL.scala 102:19]
  wire  m_1657_io_cout; // @[MUL.scala 102:19]
  wire  m_1658_io_in_0; // @[MUL.scala 124:19]
  wire  m_1658_io_in_1; // @[MUL.scala 124:19]
  wire  m_1658_io_out_0; // @[MUL.scala 124:19]
  wire  m_1658_io_out_1; // @[MUL.scala 124:19]
  wire  m_1659_io_x1; // @[MUL.scala 102:19]
  wire  m_1659_io_x2; // @[MUL.scala 102:19]
  wire  m_1659_io_x3; // @[MUL.scala 102:19]
  wire  m_1659_io_s; // @[MUL.scala 102:19]
  wire  m_1659_io_cout; // @[MUL.scala 102:19]
  wire  m_1660_io_x1; // @[MUL.scala 102:19]
  wire  m_1660_io_x2; // @[MUL.scala 102:19]
  wire  m_1660_io_x3; // @[MUL.scala 102:19]
  wire  m_1660_io_s; // @[MUL.scala 102:19]
  wire  m_1660_io_cout; // @[MUL.scala 102:19]
  wire  m_1661_io_x1; // @[MUL.scala 102:19]
  wire  m_1661_io_x2; // @[MUL.scala 102:19]
  wire  m_1661_io_x3; // @[MUL.scala 102:19]
  wire  m_1661_io_s; // @[MUL.scala 102:19]
  wire  m_1661_io_cout; // @[MUL.scala 102:19]
  wire  m_1662_io_x1; // @[MUL.scala 102:19]
  wire  m_1662_io_x2; // @[MUL.scala 102:19]
  wire  m_1662_io_x3; // @[MUL.scala 102:19]
  wire  m_1662_io_s; // @[MUL.scala 102:19]
  wire  m_1662_io_cout; // @[MUL.scala 102:19]
  wire  m_1663_io_x1; // @[MUL.scala 102:19]
  wire  m_1663_io_x2; // @[MUL.scala 102:19]
  wire  m_1663_io_x3; // @[MUL.scala 102:19]
  wire  m_1663_io_s; // @[MUL.scala 102:19]
  wire  m_1663_io_cout; // @[MUL.scala 102:19]
  wire  m_1664_io_x1; // @[MUL.scala 102:19]
  wire  m_1664_io_x2; // @[MUL.scala 102:19]
  wire  m_1664_io_x3; // @[MUL.scala 102:19]
  wire  m_1664_io_s; // @[MUL.scala 102:19]
  wire  m_1664_io_cout; // @[MUL.scala 102:19]
  wire  m_1665_io_x1; // @[MUL.scala 102:19]
  wire  m_1665_io_x2; // @[MUL.scala 102:19]
  wire  m_1665_io_x3; // @[MUL.scala 102:19]
  wire  m_1665_io_s; // @[MUL.scala 102:19]
  wire  m_1665_io_cout; // @[MUL.scala 102:19]
  wire  m_1666_io_x1; // @[MUL.scala 102:19]
  wire  m_1666_io_x2; // @[MUL.scala 102:19]
  wire  m_1666_io_x3; // @[MUL.scala 102:19]
  wire  m_1666_io_s; // @[MUL.scala 102:19]
  wire  m_1666_io_cout; // @[MUL.scala 102:19]
  wire  m_1667_io_x1; // @[MUL.scala 102:19]
  wire  m_1667_io_x2; // @[MUL.scala 102:19]
  wire  m_1667_io_x3; // @[MUL.scala 102:19]
  wire  m_1667_io_s; // @[MUL.scala 102:19]
  wire  m_1667_io_cout; // @[MUL.scala 102:19]
  wire  m_1668_io_x1; // @[MUL.scala 102:19]
  wire  m_1668_io_x2; // @[MUL.scala 102:19]
  wire  m_1668_io_x3; // @[MUL.scala 102:19]
  wire  m_1668_io_s; // @[MUL.scala 102:19]
  wire  m_1668_io_cout; // @[MUL.scala 102:19]
  wire  m_1669_io_x1; // @[MUL.scala 102:19]
  wire  m_1669_io_x2; // @[MUL.scala 102:19]
  wire  m_1669_io_x3; // @[MUL.scala 102:19]
  wire  m_1669_io_s; // @[MUL.scala 102:19]
  wire  m_1669_io_cout; // @[MUL.scala 102:19]
  wire  m_1670_io_x1; // @[MUL.scala 102:19]
  wire  m_1670_io_x2; // @[MUL.scala 102:19]
  wire  m_1670_io_x3; // @[MUL.scala 102:19]
  wire  m_1670_io_s; // @[MUL.scala 102:19]
  wire  m_1670_io_cout; // @[MUL.scala 102:19]
  wire  m_1671_io_x1; // @[MUL.scala 102:19]
  wire  m_1671_io_x2; // @[MUL.scala 102:19]
  wire  m_1671_io_x3; // @[MUL.scala 102:19]
  wire  m_1671_io_s; // @[MUL.scala 102:19]
  wire  m_1671_io_cout; // @[MUL.scala 102:19]
  wire  m_1672_io_x1; // @[MUL.scala 102:19]
  wire  m_1672_io_x2; // @[MUL.scala 102:19]
  wire  m_1672_io_x3; // @[MUL.scala 102:19]
  wire  m_1672_io_s; // @[MUL.scala 102:19]
  wire  m_1672_io_cout; // @[MUL.scala 102:19]
  wire  m_1673_io_x1; // @[MUL.scala 102:19]
  wire  m_1673_io_x2; // @[MUL.scala 102:19]
  wire  m_1673_io_x3; // @[MUL.scala 102:19]
  wire  m_1673_io_s; // @[MUL.scala 102:19]
  wire  m_1673_io_cout; // @[MUL.scala 102:19]
  wire  m_1674_io_x1; // @[MUL.scala 102:19]
  wire  m_1674_io_x2; // @[MUL.scala 102:19]
  wire  m_1674_io_x3; // @[MUL.scala 102:19]
  wire  m_1674_io_s; // @[MUL.scala 102:19]
  wire  m_1674_io_cout; // @[MUL.scala 102:19]
  wire  m_1675_io_x1; // @[MUL.scala 102:19]
  wire  m_1675_io_x2; // @[MUL.scala 102:19]
  wire  m_1675_io_x3; // @[MUL.scala 102:19]
  wire  m_1675_io_s; // @[MUL.scala 102:19]
  wire  m_1675_io_cout; // @[MUL.scala 102:19]
  wire  m_1676_io_x1; // @[MUL.scala 102:19]
  wire  m_1676_io_x2; // @[MUL.scala 102:19]
  wire  m_1676_io_x3; // @[MUL.scala 102:19]
  wire  m_1676_io_s; // @[MUL.scala 102:19]
  wire  m_1676_io_cout; // @[MUL.scala 102:19]
  wire  m_1677_io_x1; // @[MUL.scala 102:19]
  wire  m_1677_io_x2; // @[MUL.scala 102:19]
  wire  m_1677_io_x3; // @[MUL.scala 102:19]
  wire  m_1677_io_s; // @[MUL.scala 102:19]
  wire  m_1677_io_cout; // @[MUL.scala 102:19]
  wire  m_1678_io_x1; // @[MUL.scala 102:19]
  wire  m_1678_io_x2; // @[MUL.scala 102:19]
  wire  m_1678_io_x3; // @[MUL.scala 102:19]
  wire  m_1678_io_s; // @[MUL.scala 102:19]
  wire  m_1678_io_cout; // @[MUL.scala 102:19]
  wire  m_1679_io_x1; // @[MUL.scala 102:19]
  wire  m_1679_io_x2; // @[MUL.scala 102:19]
  wire  m_1679_io_x3; // @[MUL.scala 102:19]
  wire  m_1679_io_s; // @[MUL.scala 102:19]
  wire  m_1679_io_cout; // @[MUL.scala 102:19]
  wire  m_1680_io_x1; // @[MUL.scala 102:19]
  wire  m_1680_io_x2; // @[MUL.scala 102:19]
  wire  m_1680_io_x3; // @[MUL.scala 102:19]
  wire  m_1680_io_s; // @[MUL.scala 102:19]
  wire  m_1680_io_cout; // @[MUL.scala 102:19]
  wire  m_1681_io_x1; // @[MUL.scala 102:19]
  wire  m_1681_io_x2; // @[MUL.scala 102:19]
  wire  m_1681_io_x3; // @[MUL.scala 102:19]
  wire  m_1681_io_s; // @[MUL.scala 102:19]
  wire  m_1681_io_cout; // @[MUL.scala 102:19]
  wire  m_1682_io_x1; // @[MUL.scala 102:19]
  wire  m_1682_io_x2; // @[MUL.scala 102:19]
  wire  m_1682_io_x3; // @[MUL.scala 102:19]
  wire  m_1682_io_s; // @[MUL.scala 102:19]
  wire  m_1682_io_cout; // @[MUL.scala 102:19]
  wire  m_1683_io_x1; // @[MUL.scala 102:19]
  wire  m_1683_io_x2; // @[MUL.scala 102:19]
  wire  m_1683_io_x3; // @[MUL.scala 102:19]
  wire  m_1683_io_s; // @[MUL.scala 102:19]
  wire  m_1683_io_cout; // @[MUL.scala 102:19]
  wire  m_1684_io_x1; // @[MUL.scala 102:19]
  wire  m_1684_io_x2; // @[MUL.scala 102:19]
  wire  m_1684_io_x3; // @[MUL.scala 102:19]
  wire  m_1684_io_s; // @[MUL.scala 102:19]
  wire  m_1684_io_cout; // @[MUL.scala 102:19]
  wire  m_1685_io_x1; // @[MUL.scala 102:19]
  wire  m_1685_io_x2; // @[MUL.scala 102:19]
  wire  m_1685_io_x3; // @[MUL.scala 102:19]
  wire  m_1685_io_s; // @[MUL.scala 102:19]
  wire  m_1685_io_cout; // @[MUL.scala 102:19]
  wire  m_1686_io_x1; // @[MUL.scala 102:19]
  wire  m_1686_io_x2; // @[MUL.scala 102:19]
  wire  m_1686_io_x3; // @[MUL.scala 102:19]
  wire  m_1686_io_s; // @[MUL.scala 102:19]
  wire  m_1686_io_cout; // @[MUL.scala 102:19]
  wire  m_1687_io_x1; // @[MUL.scala 102:19]
  wire  m_1687_io_x2; // @[MUL.scala 102:19]
  wire  m_1687_io_x3; // @[MUL.scala 102:19]
  wire  m_1687_io_s; // @[MUL.scala 102:19]
  wire  m_1687_io_cout; // @[MUL.scala 102:19]
  wire  m_1688_io_x1; // @[MUL.scala 102:19]
  wire  m_1688_io_x2; // @[MUL.scala 102:19]
  wire  m_1688_io_x3; // @[MUL.scala 102:19]
  wire  m_1688_io_s; // @[MUL.scala 102:19]
  wire  m_1688_io_cout; // @[MUL.scala 102:19]
  wire  m_1689_io_x1; // @[MUL.scala 102:19]
  wire  m_1689_io_x2; // @[MUL.scala 102:19]
  wire  m_1689_io_x3; // @[MUL.scala 102:19]
  wire  m_1689_io_s; // @[MUL.scala 102:19]
  wire  m_1689_io_cout; // @[MUL.scala 102:19]
  wire  m_1690_io_x1; // @[MUL.scala 102:19]
  wire  m_1690_io_x2; // @[MUL.scala 102:19]
  wire  m_1690_io_x3; // @[MUL.scala 102:19]
  wire  m_1690_io_s; // @[MUL.scala 102:19]
  wire  m_1690_io_cout; // @[MUL.scala 102:19]
  wire  m_1691_io_x1; // @[MUL.scala 102:19]
  wire  m_1691_io_x2; // @[MUL.scala 102:19]
  wire  m_1691_io_x3; // @[MUL.scala 102:19]
  wire  m_1691_io_s; // @[MUL.scala 102:19]
  wire  m_1691_io_cout; // @[MUL.scala 102:19]
  wire  m_1692_io_in_0; // @[MUL.scala 124:19]
  wire  m_1692_io_in_1; // @[MUL.scala 124:19]
  wire  m_1692_io_out_0; // @[MUL.scala 124:19]
  wire  m_1692_io_out_1; // @[MUL.scala 124:19]
  wire  m_1693_io_in_0; // @[MUL.scala 124:19]
  wire  m_1693_io_in_1; // @[MUL.scala 124:19]
  wire  m_1693_io_out_0; // @[MUL.scala 124:19]
  wire  m_1693_io_out_1; // @[MUL.scala 124:19]
  wire  m_1694_io_in_0; // @[MUL.scala 124:19]
  wire  m_1694_io_in_1; // @[MUL.scala 124:19]
  wire  m_1694_io_out_0; // @[MUL.scala 124:19]
  wire  m_1694_io_out_1; // @[MUL.scala 124:19]
  wire  m_1695_io_in_0; // @[MUL.scala 124:19]
  wire  m_1695_io_in_1; // @[MUL.scala 124:19]
  wire  m_1695_io_out_0; // @[MUL.scala 124:19]
  wire  m_1695_io_out_1; // @[MUL.scala 124:19]
  wire  m_1696_io_in_0; // @[MUL.scala 124:19]
  wire  m_1696_io_in_1; // @[MUL.scala 124:19]
  wire  m_1696_io_out_0; // @[MUL.scala 124:19]
  wire  m_1696_io_out_1; // @[MUL.scala 124:19]
  wire  m_1697_io_in_0; // @[MUL.scala 124:19]
  wire  m_1697_io_in_1; // @[MUL.scala 124:19]
  wire  m_1697_io_out_0; // @[MUL.scala 124:19]
  wire  m_1697_io_out_1; // @[MUL.scala 124:19]
  wire  m_1698_io_in_0; // @[MUL.scala 124:19]
  wire  m_1698_io_in_1; // @[MUL.scala 124:19]
  wire  m_1698_io_out_0; // @[MUL.scala 124:19]
  wire  m_1698_io_out_1; // @[MUL.scala 124:19]
  wire  m_1699_io_in_0; // @[MUL.scala 124:19]
  wire  m_1699_io_in_1; // @[MUL.scala 124:19]
  wire  m_1699_io_out_0; // @[MUL.scala 124:19]
  wire  m_1699_io_out_1; // @[MUL.scala 124:19]
  wire  m_1700_io_in_0; // @[MUL.scala 124:19]
  wire  m_1700_io_in_1; // @[MUL.scala 124:19]
  wire  m_1700_io_out_0; // @[MUL.scala 124:19]
  wire  m_1700_io_out_1; // @[MUL.scala 124:19]
  wire  m_1701_io_in_0; // @[MUL.scala 124:19]
  wire  m_1701_io_in_1; // @[MUL.scala 124:19]
  wire  m_1701_io_out_0; // @[MUL.scala 124:19]
  wire  m_1701_io_out_1; // @[MUL.scala 124:19]
  wire  m_1702_io_in_0; // @[MUL.scala 124:19]
  wire  m_1702_io_in_1; // @[MUL.scala 124:19]
  wire  m_1702_io_out_0; // @[MUL.scala 124:19]
  wire  m_1702_io_out_1; // @[MUL.scala 124:19]
  wire  m_1703_io_in_0; // @[MUL.scala 124:19]
  wire  m_1703_io_in_1; // @[MUL.scala 124:19]
  wire  m_1703_io_out_0; // @[MUL.scala 124:19]
  wire  m_1703_io_out_1; // @[MUL.scala 124:19]
  wire  m_1704_io_in_0; // @[MUL.scala 124:19]
  wire  m_1704_io_in_1; // @[MUL.scala 124:19]
  wire  m_1704_io_out_0; // @[MUL.scala 124:19]
  wire  m_1704_io_out_1; // @[MUL.scala 124:19]
  wire  m_1705_io_in_0; // @[MUL.scala 124:19]
  wire  m_1705_io_in_1; // @[MUL.scala 124:19]
  wire  m_1705_io_out_0; // @[MUL.scala 124:19]
  wire  m_1705_io_out_1; // @[MUL.scala 124:19]
  wire  m_1706_io_x1; // @[MUL.scala 102:19]
  wire  m_1706_io_x2; // @[MUL.scala 102:19]
  wire  m_1706_io_x3; // @[MUL.scala 102:19]
  wire  m_1706_io_s; // @[MUL.scala 102:19]
  wire  m_1706_io_cout; // @[MUL.scala 102:19]
  wire  m_1707_io_x1; // @[MUL.scala 102:19]
  wire  m_1707_io_x2; // @[MUL.scala 102:19]
  wire  m_1707_io_x3; // @[MUL.scala 102:19]
  wire  m_1707_io_s; // @[MUL.scala 102:19]
  wire  m_1707_io_cout; // @[MUL.scala 102:19]
  wire  m_1708_io_x1; // @[MUL.scala 102:19]
  wire  m_1708_io_x2; // @[MUL.scala 102:19]
  wire  m_1708_io_x3; // @[MUL.scala 102:19]
  wire  m_1708_io_s; // @[MUL.scala 102:19]
  wire  m_1708_io_cout; // @[MUL.scala 102:19]
  wire  m_1709_io_x1; // @[MUL.scala 102:19]
  wire  m_1709_io_x2; // @[MUL.scala 102:19]
  wire  m_1709_io_x3; // @[MUL.scala 102:19]
  wire  m_1709_io_s; // @[MUL.scala 102:19]
  wire  m_1709_io_cout; // @[MUL.scala 102:19]
  wire  m_1710_io_x1; // @[MUL.scala 102:19]
  wire  m_1710_io_x2; // @[MUL.scala 102:19]
  wire  m_1710_io_x3; // @[MUL.scala 102:19]
  wire  m_1710_io_s; // @[MUL.scala 102:19]
  wire  m_1710_io_cout; // @[MUL.scala 102:19]
  wire  m_1711_io_x1; // @[MUL.scala 102:19]
  wire  m_1711_io_x2; // @[MUL.scala 102:19]
  wire  m_1711_io_x3; // @[MUL.scala 102:19]
  wire  m_1711_io_s; // @[MUL.scala 102:19]
  wire  m_1711_io_cout; // @[MUL.scala 102:19]
  wire  m_1712_io_x1; // @[MUL.scala 102:19]
  wire  m_1712_io_x2; // @[MUL.scala 102:19]
  wire  m_1712_io_x3; // @[MUL.scala 102:19]
  wire  m_1712_io_s; // @[MUL.scala 102:19]
  wire  m_1712_io_cout; // @[MUL.scala 102:19]
  wire  m_1713_io_x1; // @[MUL.scala 102:19]
  wire  m_1713_io_x2; // @[MUL.scala 102:19]
  wire  m_1713_io_x3; // @[MUL.scala 102:19]
  wire  m_1713_io_s; // @[MUL.scala 102:19]
  wire  m_1713_io_cout; // @[MUL.scala 102:19]
  wire  m_1714_io_x1; // @[MUL.scala 102:19]
  wire  m_1714_io_x2; // @[MUL.scala 102:19]
  wire  m_1714_io_x3; // @[MUL.scala 102:19]
  wire  m_1714_io_s; // @[MUL.scala 102:19]
  wire  m_1714_io_cout; // @[MUL.scala 102:19]
  wire  m_1715_io_x1; // @[MUL.scala 102:19]
  wire  m_1715_io_x2; // @[MUL.scala 102:19]
  wire  m_1715_io_x3; // @[MUL.scala 102:19]
  wire  m_1715_io_s; // @[MUL.scala 102:19]
  wire  m_1715_io_cout; // @[MUL.scala 102:19]
  wire  m_1716_io_x1; // @[MUL.scala 102:19]
  wire  m_1716_io_x2; // @[MUL.scala 102:19]
  wire  m_1716_io_x3; // @[MUL.scala 102:19]
  wire  m_1716_io_s; // @[MUL.scala 102:19]
  wire  m_1716_io_cout; // @[MUL.scala 102:19]
  wire  m_1717_io_x1; // @[MUL.scala 102:19]
  wire  m_1717_io_x2; // @[MUL.scala 102:19]
  wire  m_1717_io_x3; // @[MUL.scala 102:19]
  wire  m_1717_io_s; // @[MUL.scala 102:19]
  wire  m_1717_io_cout; // @[MUL.scala 102:19]
  wire  m_1718_io_x1; // @[MUL.scala 102:19]
  wire  m_1718_io_x2; // @[MUL.scala 102:19]
  wire  m_1718_io_x3; // @[MUL.scala 102:19]
  wire  m_1718_io_s; // @[MUL.scala 102:19]
  wire  m_1718_io_cout; // @[MUL.scala 102:19]
  wire  m_1719_io_x1; // @[MUL.scala 102:19]
  wire  m_1719_io_x2; // @[MUL.scala 102:19]
  wire  m_1719_io_x3; // @[MUL.scala 102:19]
  wire  m_1719_io_s; // @[MUL.scala 102:19]
  wire  m_1719_io_cout; // @[MUL.scala 102:19]
  wire  m_1720_io_x1; // @[MUL.scala 102:19]
  wire  m_1720_io_x2; // @[MUL.scala 102:19]
  wire  m_1720_io_x3; // @[MUL.scala 102:19]
  wire  m_1720_io_s; // @[MUL.scala 102:19]
  wire  m_1720_io_cout; // @[MUL.scala 102:19]
  wire  m_1721_io_in_0; // @[MUL.scala 124:19]
  wire  m_1721_io_in_1; // @[MUL.scala 124:19]
  wire  m_1721_io_out_0; // @[MUL.scala 124:19]
  wire  m_1721_io_out_1; // @[MUL.scala 124:19]
  wire  m_1722_io_x1; // @[MUL.scala 102:19]
  wire  m_1722_io_x2; // @[MUL.scala 102:19]
  wire  m_1722_io_x3; // @[MUL.scala 102:19]
  wire  m_1722_io_s; // @[MUL.scala 102:19]
  wire  m_1722_io_cout; // @[MUL.scala 102:19]
  wire  m_1723_io_in_0; // @[MUL.scala 124:19]
  wire  m_1723_io_in_1; // @[MUL.scala 124:19]
  wire  m_1723_io_out_0; // @[MUL.scala 124:19]
  wire  m_1723_io_out_1; // @[MUL.scala 124:19]
  wire  m_1724_io_x1; // @[MUL.scala 102:19]
  wire  m_1724_io_x2; // @[MUL.scala 102:19]
  wire  m_1724_io_x3; // @[MUL.scala 102:19]
  wire  m_1724_io_s; // @[MUL.scala 102:19]
  wire  m_1724_io_cout; // @[MUL.scala 102:19]
  wire  m_1725_io_in_0; // @[MUL.scala 124:19]
  wire  m_1725_io_in_1; // @[MUL.scala 124:19]
  wire  m_1725_io_out_0; // @[MUL.scala 124:19]
  wire  m_1725_io_out_1; // @[MUL.scala 124:19]
  wire  m_1726_io_x1; // @[MUL.scala 102:19]
  wire  m_1726_io_x2; // @[MUL.scala 102:19]
  wire  m_1726_io_x3; // @[MUL.scala 102:19]
  wire  m_1726_io_s; // @[MUL.scala 102:19]
  wire  m_1726_io_cout; // @[MUL.scala 102:19]
  wire  m_1727_io_in_0; // @[MUL.scala 124:19]
  wire  m_1727_io_in_1; // @[MUL.scala 124:19]
  wire  m_1727_io_out_0; // @[MUL.scala 124:19]
  wire  m_1727_io_out_1; // @[MUL.scala 124:19]
  wire  m_1728_io_x1; // @[MUL.scala 102:19]
  wire  m_1728_io_x2; // @[MUL.scala 102:19]
  wire  m_1728_io_x3; // @[MUL.scala 102:19]
  wire  m_1728_io_s; // @[MUL.scala 102:19]
  wire  m_1728_io_cout; // @[MUL.scala 102:19]
  wire  m_1729_io_in_0; // @[MUL.scala 124:19]
  wire  m_1729_io_in_1; // @[MUL.scala 124:19]
  wire  m_1729_io_out_0; // @[MUL.scala 124:19]
  wire  m_1729_io_out_1; // @[MUL.scala 124:19]
  wire  m_1730_io_x1; // @[MUL.scala 102:19]
  wire  m_1730_io_x2; // @[MUL.scala 102:19]
  wire  m_1730_io_x3; // @[MUL.scala 102:19]
  wire  m_1730_io_s; // @[MUL.scala 102:19]
  wire  m_1730_io_cout; // @[MUL.scala 102:19]
  wire  m_1731_io_x1; // @[MUL.scala 102:19]
  wire  m_1731_io_x2; // @[MUL.scala 102:19]
  wire  m_1731_io_x3; // @[MUL.scala 102:19]
  wire  m_1731_io_s; // @[MUL.scala 102:19]
  wire  m_1731_io_cout; // @[MUL.scala 102:19]
  wire  m_1732_io_x1; // @[MUL.scala 102:19]
  wire  m_1732_io_x2; // @[MUL.scala 102:19]
  wire  m_1732_io_x3; // @[MUL.scala 102:19]
  wire  m_1732_io_s; // @[MUL.scala 102:19]
  wire  m_1732_io_cout; // @[MUL.scala 102:19]
  wire  m_1733_io_x1; // @[MUL.scala 102:19]
  wire  m_1733_io_x2; // @[MUL.scala 102:19]
  wire  m_1733_io_x3; // @[MUL.scala 102:19]
  wire  m_1733_io_s; // @[MUL.scala 102:19]
  wire  m_1733_io_cout; // @[MUL.scala 102:19]
  wire  m_1734_io_x1; // @[MUL.scala 102:19]
  wire  m_1734_io_x2; // @[MUL.scala 102:19]
  wire  m_1734_io_x3; // @[MUL.scala 102:19]
  wire  m_1734_io_s; // @[MUL.scala 102:19]
  wire  m_1734_io_cout; // @[MUL.scala 102:19]
  wire  m_1735_io_x1; // @[MUL.scala 102:19]
  wire  m_1735_io_x2; // @[MUL.scala 102:19]
  wire  m_1735_io_x3; // @[MUL.scala 102:19]
  wire  m_1735_io_s; // @[MUL.scala 102:19]
  wire  m_1735_io_cout; // @[MUL.scala 102:19]
  wire  m_1736_io_x1; // @[MUL.scala 102:19]
  wire  m_1736_io_x2; // @[MUL.scala 102:19]
  wire  m_1736_io_x3; // @[MUL.scala 102:19]
  wire  m_1736_io_s; // @[MUL.scala 102:19]
  wire  m_1736_io_cout; // @[MUL.scala 102:19]
  wire  m_1737_io_x1; // @[MUL.scala 102:19]
  wire  m_1737_io_x2; // @[MUL.scala 102:19]
  wire  m_1737_io_x3; // @[MUL.scala 102:19]
  wire  m_1737_io_s; // @[MUL.scala 102:19]
  wire  m_1737_io_cout; // @[MUL.scala 102:19]
  wire  m_1738_io_x1; // @[MUL.scala 102:19]
  wire  m_1738_io_x2; // @[MUL.scala 102:19]
  wire  m_1738_io_x3; // @[MUL.scala 102:19]
  wire  m_1738_io_s; // @[MUL.scala 102:19]
  wire  m_1738_io_cout; // @[MUL.scala 102:19]
  wire  m_1739_io_x1; // @[MUL.scala 102:19]
  wire  m_1739_io_x2; // @[MUL.scala 102:19]
  wire  m_1739_io_x3; // @[MUL.scala 102:19]
  wire  m_1739_io_s; // @[MUL.scala 102:19]
  wire  m_1739_io_cout; // @[MUL.scala 102:19]
  wire  m_1740_io_x1; // @[MUL.scala 102:19]
  wire  m_1740_io_x2; // @[MUL.scala 102:19]
  wire  m_1740_io_x3; // @[MUL.scala 102:19]
  wire  m_1740_io_s; // @[MUL.scala 102:19]
  wire  m_1740_io_cout; // @[MUL.scala 102:19]
  wire  m_1741_io_x1; // @[MUL.scala 102:19]
  wire  m_1741_io_x2; // @[MUL.scala 102:19]
  wire  m_1741_io_x3; // @[MUL.scala 102:19]
  wire  m_1741_io_s; // @[MUL.scala 102:19]
  wire  m_1741_io_cout; // @[MUL.scala 102:19]
  wire  m_1742_io_x1; // @[MUL.scala 102:19]
  wire  m_1742_io_x2; // @[MUL.scala 102:19]
  wire  m_1742_io_x3; // @[MUL.scala 102:19]
  wire  m_1742_io_s; // @[MUL.scala 102:19]
  wire  m_1742_io_cout; // @[MUL.scala 102:19]
  wire  m_1743_io_x1; // @[MUL.scala 102:19]
  wire  m_1743_io_x2; // @[MUL.scala 102:19]
  wire  m_1743_io_x3; // @[MUL.scala 102:19]
  wire  m_1743_io_s; // @[MUL.scala 102:19]
  wire  m_1743_io_cout; // @[MUL.scala 102:19]
  wire  m_1744_io_x1; // @[MUL.scala 102:19]
  wire  m_1744_io_x2; // @[MUL.scala 102:19]
  wire  m_1744_io_x3; // @[MUL.scala 102:19]
  wire  m_1744_io_s; // @[MUL.scala 102:19]
  wire  m_1744_io_cout; // @[MUL.scala 102:19]
  wire  m_1745_io_x1; // @[MUL.scala 102:19]
  wire  m_1745_io_x2; // @[MUL.scala 102:19]
  wire  m_1745_io_x3; // @[MUL.scala 102:19]
  wire  m_1745_io_s; // @[MUL.scala 102:19]
  wire  m_1745_io_cout; // @[MUL.scala 102:19]
  wire  m_1746_io_x1; // @[MUL.scala 102:19]
  wire  m_1746_io_x2; // @[MUL.scala 102:19]
  wire  m_1746_io_x3; // @[MUL.scala 102:19]
  wire  m_1746_io_s; // @[MUL.scala 102:19]
  wire  m_1746_io_cout; // @[MUL.scala 102:19]
  wire  m_1747_io_x1; // @[MUL.scala 102:19]
  wire  m_1747_io_x2; // @[MUL.scala 102:19]
  wire  m_1747_io_x3; // @[MUL.scala 102:19]
  wire  m_1747_io_s; // @[MUL.scala 102:19]
  wire  m_1747_io_cout; // @[MUL.scala 102:19]
  wire  m_1748_io_x1; // @[MUL.scala 102:19]
  wire  m_1748_io_x2; // @[MUL.scala 102:19]
  wire  m_1748_io_x3; // @[MUL.scala 102:19]
  wire  m_1748_io_s; // @[MUL.scala 102:19]
  wire  m_1748_io_cout; // @[MUL.scala 102:19]
  wire  m_1749_io_x1; // @[MUL.scala 102:19]
  wire  m_1749_io_x2; // @[MUL.scala 102:19]
  wire  m_1749_io_x3; // @[MUL.scala 102:19]
  wire  m_1749_io_s; // @[MUL.scala 102:19]
  wire  m_1749_io_cout; // @[MUL.scala 102:19]
  wire  m_1750_io_x1; // @[MUL.scala 102:19]
  wire  m_1750_io_x2; // @[MUL.scala 102:19]
  wire  m_1750_io_x3; // @[MUL.scala 102:19]
  wire  m_1750_io_s; // @[MUL.scala 102:19]
  wire  m_1750_io_cout; // @[MUL.scala 102:19]
  wire  m_1751_io_x1; // @[MUL.scala 102:19]
  wire  m_1751_io_x2; // @[MUL.scala 102:19]
  wire  m_1751_io_x3; // @[MUL.scala 102:19]
  wire  m_1751_io_s; // @[MUL.scala 102:19]
  wire  m_1751_io_cout; // @[MUL.scala 102:19]
  wire  m_1752_io_x1; // @[MUL.scala 102:19]
  wire  m_1752_io_x2; // @[MUL.scala 102:19]
  wire  m_1752_io_x3; // @[MUL.scala 102:19]
  wire  m_1752_io_s; // @[MUL.scala 102:19]
  wire  m_1752_io_cout; // @[MUL.scala 102:19]
  wire  m_1753_io_x1; // @[MUL.scala 102:19]
  wire  m_1753_io_x2; // @[MUL.scala 102:19]
  wire  m_1753_io_x3; // @[MUL.scala 102:19]
  wire  m_1753_io_s; // @[MUL.scala 102:19]
  wire  m_1753_io_cout; // @[MUL.scala 102:19]
  wire  m_1754_io_x1; // @[MUL.scala 102:19]
  wire  m_1754_io_x2; // @[MUL.scala 102:19]
  wire  m_1754_io_x3; // @[MUL.scala 102:19]
  wire  m_1754_io_s; // @[MUL.scala 102:19]
  wire  m_1754_io_cout; // @[MUL.scala 102:19]
  wire  m_1755_io_x1; // @[MUL.scala 102:19]
  wire  m_1755_io_x2; // @[MUL.scala 102:19]
  wire  m_1755_io_x3; // @[MUL.scala 102:19]
  wire  m_1755_io_s; // @[MUL.scala 102:19]
  wire  m_1755_io_cout; // @[MUL.scala 102:19]
  wire  m_1756_io_x1; // @[MUL.scala 102:19]
  wire  m_1756_io_x2; // @[MUL.scala 102:19]
  wire  m_1756_io_x3; // @[MUL.scala 102:19]
  wire  m_1756_io_s; // @[MUL.scala 102:19]
  wire  m_1756_io_cout; // @[MUL.scala 102:19]
  wire  m_1757_io_x1; // @[MUL.scala 102:19]
  wire  m_1757_io_x2; // @[MUL.scala 102:19]
  wire  m_1757_io_x3; // @[MUL.scala 102:19]
  wire  m_1757_io_s; // @[MUL.scala 102:19]
  wire  m_1757_io_cout; // @[MUL.scala 102:19]
  wire  m_1758_io_x1; // @[MUL.scala 102:19]
  wire  m_1758_io_x2; // @[MUL.scala 102:19]
  wire  m_1758_io_x3; // @[MUL.scala 102:19]
  wire  m_1758_io_s; // @[MUL.scala 102:19]
  wire  m_1758_io_cout; // @[MUL.scala 102:19]
  wire  m_1759_io_x1; // @[MUL.scala 102:19]
  wire  m_1759_io_x2; // @[MUL.scala 102:19]
  wire  m_1759_io_x3; // @[MUL.scala 102:19]
  wire  m_1759_io_s; // @[MUL.scala 102:19]
  wire  m_1759_io_cout; // @[MUL.scala 102:19]
  wire  m_1760_io_in_0; // @[MUL.scala 124:19]
  wire  m_1760_io_in_1; // @[MUL.scala 124:19]
  wire  m_1760_io_out_0; // @[MUL.scala 124:19]
  wire  m_1760_io_out_1; // @[MUL.scala 124:19]
  wire  m_1761_io_x1; // @[MUL.scala 102:19]
  wire  m_1761_io_x2; // @[MUL.scala 102:19]
  wire  m_1761_io_x3; // @[MUL.scala 102:19]
  wire  m_1761_io_s; // @[MUL.scala 102:19]
  wire  m_1761_io_cout; // @[MUL.scala 102:19]
  wire  m_1762_io_x1; // @[MUL.scala 102:19]
  wire  m_1762_io_x2; // @[MUL.scala 102:19]
  wire  m_1762_io_x3; // @[MUL.scala 102:19]
  wire  m_1762_io_s; // @[MUL.scala 102:19]
  wire  m_1762_io_cout; // @[MUL.scala 102:19]
  wire  m_1763_io_in_0; // @[MUL.scala 124:19]
  wire  m_1763_io_in_1; // @[MUL.scala 124:19]
  wire  m_1763_io_out_0; // @[MUL.scala 124:19]
  wire  m_1763_io_out_1; // @[MUL.scala 124:19]
  wire  m_1764_io_x1; // @[MUL.scala 102:19]
  wire  m_1764_io_x2; // @[MUL.scala 102:19]
  wire  m_1764_io_x3; // @[MUL.scala 102:19]
  wire  m_1764_io_s; // @[MUL.scala 102:19]
  wire  m_1764_io_cout; // @[MUL.scala 102:19]
  wire  m_1765_io_x1; // @[MUL.scala 102:19]
  wire  m_1765_io_x2; // @[MUL.scala 102:19]
  wire  m_1765_io_x3; // @[MUL.scala 102:19]
  wire  m_1765_io_s; // @[MUL.scala 102:19]
  wire  m_1765_io_cout; // @[MUL.scala 102:19]
  wire  m_1766_io_in_0; // @[MUL.scala 124:19]
  wire  m_1766_io_in_1; // @[MUL.scala 124:19]
  wire  m_1766_io_out_0; // @[MUL.scala 124:19]
  wire  m_1766_io_out_1; // @[MUL.scala 124:19]
  wire  m_1767_io_x1; // @[MUL.scala 102:19]
  wire  m_1767_io_x2; // @[MUL.scala 102:19]
  wire  m_1767_io_x3; // @[MUL.scala 102:19]
  wire  m_1767_io_s; // @[MUL.scala 102:19]
  wire  m_1767_io_cout; // @[MUL.scala 102:19]
  wire  m_1768_io_x1; // @[MUL.scala 102:19]
  wire  m_1768_io_x2; // @[MUL.scala 102:19]
  wire  m_1768_io_x3; // @[MUL.scala 102:19]
  wire  m_1768_io_s; // @[MUL.scala 102:19]
  wire  m_1768_io_cout; // @[MUL.scala 102:19]
  wire  m_1769_io_in_0; // @[MUL.scala 124:19]
  wire  m_1769_io_in_1; // @[MUL.scala 124:19]
  wire  m_1769_io_out_0; // @[MUL.scala 124:19]
  wire  m_1769_io_out_1; // @[MUL.scala 124:19]
  wire  m_1770_io_x1; // @[MUL.scala 102:19]
  wire  m_1770_io_x2; // @[MUL.scala 102:19]
  wire  m_1770_io_x3; // @[MUL.scala 102:19]
  wire  m_1770_io_s; // @[MUL.scala 102:19]
  wire  m_1770_io_cout; // @[MUL.scala 102:19]
  wire  m_1771_io_x1; // @[MUL.scala 102:19]
  wire  m_1771_io_x2; // @[MUL.scala 102:19]
  wire  m_1771_io_x3; // @[MUL.scala 102:19]
  wire  m_1771_io_s; // @[MUL.scala 102:19]
  wire  m_1771_io_cout; // @[MUL.scala 102:19]
  wire  m_1772_io_in_0; // @[MUL.scala 124:19]
  wire  m_1772_io_in_1; // @[MUL.scala 124:19]
  wire  m_1772_io_out_0; // @[MUL.scala 124:19]
  wire  m_1772_io_out_1; // @[MUL.scala 124:19]
  wire  m_1773_io_x1; // @[MUL.scala 102:19]
  wire  m_1773_io_x2; // @[MUL.scala 102:19]
  wire  m_1773_io_x3; // @[MUL.scala 102:19]
  wire  m_1773_io_s; // @[MUL.scala 102:19]
  wire  m_1773_io_cout; // @[MUL.scala 102:19]
  wire  m_1774_io_x1; // @[MUL.scala 102:19]
  wire  m_1774_io_x2; // @[MUL.scala 102:19]
  wire  m_1774_io_x3; // @[MUL.scala 102:19]
  wire  m_1774_io_s; // @[MUL.scala 102:19]
  wire  m_1774_io_cout; // @[MUL.scala 102:19]
  wire  m_1775_io_in_0; // @[MUL.scala 124:19]
  wire  m_1775_io_in_1; // @[MUL.scala 124:19]
  wire  m_1775_io_out_0; // @[MUL.scala 124:19]
  wire  m_1775_io_out_1; // @[MUL.scala 124:19]
  wire  m_1776_io_x1; // @[MUL.scala 102:19]
  wire  m_1776_io_x2; // @[MUL.scala 102:19]
  wire  m_1776_io_x3; // @[MUL.scala 102:19]
  wire  m_1776_io_s; // @[MUL.scala 102:19]
  wire  m_1776_io_cout; // @[MUL.scala 102:19]
  wire  m_1777_io_x1; // @[MUL.scala 102:19]
  wire  m_1777_io_x2; // @[MUL.scala 102:19]
  wire  m_1777_io_x3; // @[MUL.scala 102:19]
  wire  m_1777_io_s; // @[MUL.scala 102:19]
  wire  m_1777_io_cout; // @[MUL.scala 102:19]
  wire  m_1778_io_in_0; // @[MUL.scala 124:19]
  wire  m_1778_io_in_1; // @[MUL.scala 124:19]
  wire  m_1778_io_out_0; // @[MUL.scala 124:19]
  wire  m_1778_io_out_1; // @[MUL.scala 124:19]
  wire  m_1779_io_x1; // @[MUL.scala 102:19]
  wire  m_1779_io_x2; // @[MUL.scala 102:19]
  wire  m_1779_io_x3; // @[MUL.scala 102:19]
  wire  m_1779_io_s; // @[MUL.scala 102:19]
  wire  m_1779_io_cout; // @[MUL.scala 102:19]
  wire  m_1780_io_x1; // @[MUL.scala 102:19]
  wire  m_1780_io_x2; // @[MUL.scala 102:19]
  wire  m_1780_io_x3; // @[MUL.scala 102:19]
  wire  m_1780_io_s; // @[MUL.scala 102:19]
  wire  m_1780_io_cout; // @[MUL.scala 102:19]
  wire  m_1781_io_in_0; // @[MUL.scala 124:19]
  wire  m_1781_io_in_1; // @[MUL.scala 124:19]
  wire  m_1781_io_out_0; // @[MUL.scala 124:19]
  wire  m_1781_io_out_1; // @[MUL.scala 124:19]
  wire  m_1782_io_x1; // @[MUL.scala 102:19]
  wire  m_1782_io_x2; // @[MUL.scala 102:19]
  wire  m_1782_io_x3; // @[MUL.scala 102:19]
  wire  m_1782_io_s; // @[MUL.scala 102:19]
  wire  m_1782_io_cout; // @[MUL.scala 102:19]
  wire  m_1783_io_x1; // @[MUL.scala 102:19]
  wire  m_1783_io_x2; // @[MUL.scala 102:19]
  wire  m_1783_io_x3; // @[MUL.scala 102:19]
  wire  m_1783_io_s; // @[MUL.scala 102:19]
  wire  m_1783_io_cout; // @[MUL.scala 102:19]
  wire  m_1784_io_x1; // @[MUL.scala 102:19]
  wire  m_1784_io_x2; // @[MUL.scala 102:19]
  wire  m_1784_io_x3; // @[MUL.scala 102:19]
  wire  m_1784_io_s; // @[MUL.scala 102:19]
  wire  m_1784_io_cout; // @[MUL.scala 102:19]
  wire  m_1785_io_x1; // @[MUL.scala 102:19]
  wire  m_1785_io_x2; // @[MUL.scala 102:19]
  wire  m_1785_io_x3; // @[MUL.scala 102:19]
  wire  m_1785_io_s; // @[MUL.scala 102:19]
  wire  m_1785_io_cout; // @[MUL.scala 102:19]
  wire  m_1786_io_x1; // @[MUL.scala 102:19]
  wire  m_1786_io_x2; // @[MUL.scala 102:19]
  wire  m_1786_io_x3; // @[MUL.scala 102:19]
  wire  m_1786_io_s; // @[MUL.scala 102:19]
  wire  m_1786_io_cout; // @[MUL.scala 102:19]
  wire  m_1787_io_x1; // @[MUL.scala 102:19]
  wire  m_1787_io_x2; // @[MUL.scala 102:19]
  wire  m_1787_io_x3; // @[MUL.scala 102:19]
  wire  m_1787_io_s; // @[MUL.scala 102:19]
  wire  m_1787_io_cout; // @[MUL.scala 102:19]
  wire  m_1788_io_x1; // @[MUL.scala 102:19]
  wire  m_1788_io_x2; // @[MUL.scala 102:19]
  wire  m_1788_io_x3; // @[MUL.scala 102:19]
  wire  m_1788_io_s; // @[MUL.scala 102:19]
  wire  m_1788_io_cout; // @[MUL.scala 102:19]
  wire  m_1789_io_x1; // @[MUL.scala 102:19]
  wire  m_1789_io_x2; // @[MUL.scala 102:19]
  wire  m_1789_io_x3; // @[MUL.scala 102:19]
  wire  m_1789_io_s; // @[MUL.scala 102:19]
  wire  m_1789_io_cout; // @[MUL.scala 102:19]
  wire  m_1790_io_x1; // @[MUL.scala 102:19]
  wire  m_1790_io_x2; // @[MUL.scala 102:19]
  wire  m_1790_io_x3; // @[MUL.scala 102:19]
  wire  m_1790_io_s; // @[MUL.scala 102:19]
  wire  m_1790_io_cout; // @[MUL.scala 102:19]
  wire  m_1791_io_x1; // @[MUL.scala 102:19]
  wire  m_1791_io_x2; // @[MUL.scala 102:19]
  wire  m_1791_io_x3; // @[MUL.scala 102:19]
  wire  m_1791_io_s; // @[MUL.scala 102:19]
  wire  m_1791_io_cout; // @[MUL.scala 102:19]
  wire  m_1792_io_x1; // @[MUL.scala 102:19]
  wire  m_1792_io_x2; // @[MUL.scala 102:19]
  wire  m_1792_io_x3; // @[MUL.scala 102:19]
  wire  m_1792_io_s; // @[MUL.scala 102:19]
  wire  m_1792_io_cout; // @[MUL.scala 102:19]
  wire  m_1793_io_x1; // @[MUL.scala 102:19]
  wire  m_1793_io_x2; // @[MUL.scala 102:19]
  wire  m_1793_io_x3; // @[MUL.scala 102:19]
  wire  m_1793_io_s; // @[MUL.scala 102:19]
  wire  m_1793_io_cout; // @[MUL.scala 102:19]
  wire  m_1794_io_x1; // @[MUL.scala 102:19]
  wire  m_1794_io_x2; // @[MUL.scala 102:19]
  wire  m_1794_io_x3; // @[MUL.scala 102:19]
  wire  m_1794_io_s; // @[MUL.scala 102:19]
  wire  m_1794_io_cout; // @[MUL.scala 102:19]
  wire  m_1795_io_x1; // @[MUL.scala 102:19]
  wire  m_1795_io_x2; // @[MUL.scala 102:19]
  wire  m_1795_io_x3; // @[MUL.scala 102:19]
  wire  m_1795_io_s; // @[MUL.scala 102:19]
  wire  m_1795_io_cout; // @[MUL.scala 102:19]
  wire  m_1796_io_x1; // @[MUL.scala 102:19]
  wire  m_1796_io_x2; // @[MUL.scala 102:19]
  wire  m_1796_io_x3; // @[MUL.scala 102:19]
  wire  m_1796_io_s; // @[MUL.scala 102:19]
  wire  m_1796_io_cout; // @[MUL.scala 102:19]
  wire  m_1797_io_x1; // @[MUL.scala 102:19]
  wire  m_1797_io_x2; // @[MUL.scala 102:19]
  wire  m_1797_io_x3; // @[MUL.scala 102:19]
  wire  m_1797_io_s; // @[MUL.scala 102:19]
  wire  m_1797_io_cout; // @[MUL.scala 102:19]
  wire  m_1798_io_x1; // @[MUL.scala 102:19]
  wire  m_1798_io_x2; // @[MUL.scala 102:19]
  wire  m_1798_io_x3; // @[MUL.scala 102:19]
  wire  m_1798_io_s; // @[MUL.scala 102:19]
  wire  m_1798_io_cout; // @[MUL.scala 102:19]
  wire  m_1799_io_x1; // @[MUL.scala 102:19]
  wire  m_1799_io_x2; // @[MUL.scala 102:19]
  wire  m_1799_io_x3; // @[MUL.scala 102:19]
  wire  m_1799_io_s; // @[MUL.scala 102:19]
  wire  m_1799_io_cout; // @[MUL.scala 102:19]
  wire  m_1800_io_x1; // @[MUL.scala 102:19]
  wire  m_1800_io_x2; // @[MUL.scala 102:19]
  wire  m_1800_io_x3; // @[MUL.scala 102:19]
  wire  m_1800_io_s; // @[MUL.scala 102:19]
  wire  m_1800_io_cout; // @[MUL.scala 102:19]
  wire  m_1801_io_x1; // @[MUL.scala 102:19]
  wire  m_1801_io_x2; // @[MUL.scala 102:19]
  wire  m_1801_io_x3; // @[MUL.scala 102:19]
  wire  m_1801_io_s; // @[MUL.scala 102:19]
  wire  m_1801_io_cout; // @[MUL.scala 102:19]
  wire  m_1802_io_x1; // @[MUL.scala 102:19]
  wire  m_1802_io_x2; // @[MUL.scala 102:19]
  wire  m_1802_io_x3; // @[MUL.scala 102:19]
  wire  m_1802_io_s; // @[MUL.scala 102:19]
  wire  m_1802_io_cout; // @[MUL.scala 102:19]
  wire  m_1803_io_x1; // @[MUL.scala 102:19]
  wire  m_1803_io_x2; // @[MUL.scala 102:19]
  wire  m_1803_io_x3; // @[MUL.scala 102:19]
  wire  m_1803_io_s; // @[MUL.scala 102:19]
  wire  m_1803_io_cout; // @[MUL.scala 102:19]
  wire  m_1804_io_x1; // @[MUL.scala 102:19]
  wire  m_1804_io_x2; // @[MUL.scala 102:19]
  wire  m_1804_io_x3; // @[MUL.scala 102:19]
  wire  m_1804_io_s; // @[MUL.scala 102:19]
  wire  m_1804_io_cout; // @[MUL.scala 102:19]
  wire  m_1805_io_x1; // @[MUL.scala 102:19]
  wire  m_1805_io_x2; // @[MUL.scala 102:19]
  wire  m_1805_io_x3; // @[MUL.scala 102:19]
  wire  m_1805_io_s; // @[MUL.scala 102:19]
  wire  m_1805_io_cout; // @[MUL.scala 102:19]
  wire  m_1806_io_x1; // @[MUL.scala 102:19]
  wire  m_1806_io_x2; // @[MUL.scala 102:19]
  wire  m_1806_io_x3; // @[MUL.scala 102:19]
  wire  m_1806_io_s; // @[MUL.scala 102:19]
  wire  m_1806_io_cout; // @[MUL.scala 102:19]
  wire  m_1807_io_x1; // @[MUL.scala 102:19]
  wire  m_1807_io_x2; // @[MUL.scala 102:19]
  wire  m_1807_io_x3; // @[MUL.scala 102:19]
  wire  m_1807_io_s; // @[MUL.scala 102:19]
  wire  m_1807_io_cout; // @[MUL.scala 102:19]
  wire  m_1808_io_x1; // @[MUL.scala 102:19]
  wire  m_1808_io_x2; // @[MUL.scala 102:19]
  wire  m_1808_io_x3; // @[MUL.scala 102:19]
  wire  m_1808_io_s; // @[MUL.scala 102:19]
  wire  m_1808_io_cout; // @[MUL.scala 102:19]
  wire  m_1809_io_x1; // @[MUL.scala 102:19]
  wire  m_1809_io_x2; // @[MUL.scala 102:19]
  wire  m_1809_io_x3; // @[MUL.scala 102:19]
  wire  m_1809_io_s; // @[MUL.scala 102:19]
  wire  m_1809_io_cout; // @[MUL.scala 102:19]
  wire  m_1810_io_x1; // @[MUL.scala 102:19]
  wire  m_1810_io_x2; // @[MUL.scala 102:19]
  wire  m_1810_io_x3; // @[MUL.scala 102:19]
  wire  m_1810_io_s; // @[MUL.scala 102:19]
  wire  m_1810_io_cout; // @[MUL.scala 102:19]
  wire  m_1811_io_x1; // @[MUL.scala 102:19]
  wire  m_1811_io_x2; // @[MUL.scala 102:19]
  wire  m_1811_io_x3; // @[MUL.scala 102:19]
  wire  m_1811_io_s; // @[MUL.scala 102:19]
  wire  m_1811_io_cout; // @[MUL.scala 102:19]
  wire  m_1812_io_x1; // @[MUL.scala 102:19]
  wire  m_1812_io_x2; // @[MUL.scala 102:19]
  wire  m_1812_io_x3; // @[MUL.scala 102:19]
  wire  m_1812_io_s; // @[MUL.scala 102:19]
  wire  m_1812_io_cout; // @[MUL.scala 102:19]
  wire  m_1813_io_x1; // @[MUL.scala 102:19]
  wire  m_1813_io_x2; // @[MUL.scala 102:19]
  wire  m_1813_io_x3; // @[MUL.scala 102:19]
  wire  m_1813_io_s; // @[MUL.scala 102:19]
  wire  m_1813_io_cout; // @[MUL.scala 102:19]
  wire  m_1814_io_x1; // @[MUL.scala 102:19]
  wire  m_1814_io_x2; // @[MUL.scala 102:19]
  wire  m_1814_io_x3; // @[MUL.scala 102:19]
  wire  m_1814_io_s; // @[MUL.scala 102:19]
  wire  m_1814_io_cout; // @[MUL.scala 102:19]
  wire  m_1815_io_x1; // @[MUL.scala 102:19]
  wire  m_1815_io_x2; // @[MUL.scala 102:19]
  wire  m_1815_io_x3; // @[MUL.scala 102:19]
  wire  m_1815_io_s; // @[MUL.scala 102:19]
  wire  m_1815_io_cout; // @[MUL.scala 102:19]
  wire  m_1816_io_x1; // @[MUL.scala 102:19]
  wire  m_1816_io_x2; // @[MUL.scala 102:19]
  wire  m_1816_io_x3; // @[MUL.scala 102:19]
  wire  m_1816_io_s; // @[MUL.scala 102:19]
  wire  m_1816_io_cout; // @[MUL.scala 102:19]
  wire  m_1817_io_x1; // @[MUL.scala 102:19]
  wire  m_1817_io_x2; // @[MUL.scala 102:19]
  wire  m_1817_io_x3; // @[MUL.scala 102:19]
  wire  m_1817_io_s; // @[MUL.scala 102:19]
  wire  m_1817_io_cout; // @[MUL.scala 102:19]
  wire  m_1818_io_x1; // @[MUL.scala 102:19]
  wire  m_1818_io_x2; // @[MUL.scala 102:19]
  wire  m_1818_io_x3; // @[MUL.scala 102:19]
  wire  m_1818_io_s; // @[MUL.scala 102:19]
  wire  m_1818_io_cout; // @[MUL.scala 102:19]
  wire  m_1819_io_x1; // @[MUL.scala 102:19]
  wire  m_1819_io_x2; // @[MUL.scala 102:19]
  wire  m_1819_io_x3; // @[MUL.scala 102:19]
  wire  m_1819_io_s; // @[MUL.scala 102:19]
  wire  m_1819_io_cout; // @[MUL.scala 102:19]
  wire  m_1820_io_x1; // @[MUL.scala 102:19]
  wire  m_1820_io_x2; // @[MUL.scala 102:19]
  wire  m_1820_io_x3; // @[MUL.scala 102:19]
  wire  m_1820_io_s; // @[MUL.scala 102:19]
  wire  m_1820_io_cout; // @[MUL.scala 102:19]
  wire  m_1821_io_x1; // @[MUL.scala 102:19]
  wire  m_1821_io_x2; // @[MUL.scala 102:19]
  wire  m_1821_io_x3; // @[MUL.scala 102:19]
  wire  m_1821_io_s; // @[MUL.scala 102:19]
  wire  m_1821_io_cout; // @[MUL.scala 102:19]
  wire  m_1822_io_x1; // @[MUL.scala 102:19]
  wire  m_1822_io_x2; // @[MUL.scala 102:19]
  wire  m_1822_io_x3; // @[MUL.scala 102:19]
  wire  m_1822_io_s; // @[MUL.scala 102:19]
  wire  m_1822_io_cout; // @[MUL.scala 102:19]
  wire  m_1823_io_x1; // @[MUL.scala 102:19]
  wire  m_1823_io_x2; // @[MUL.scala 102:19]
  wire  m_1823_io_x3; // @[MUL.scala 102:19]
  wire  m_1823_io_s; // @[MUL.scala 102:19]
  wire  m_1823_io_cout; // @[MUL.scala 102:19]
  wire  m_1824_io_x1; // @[MUL.scala 102:19]
  wire  m_1824_io_x2; // @[MUL.scala 102:19]
  wire  m_1824_io_x3; // @[MUL.scala 102:19]
  wire  m_1824_io_s; // @[MUL.scala 102:19]
  wire  m_1824_io_cout; // @[MUL.scala 102:19]
  wire  m_1825_io_x1; // @[MUL.scala 102:19]
  wire  m_1825_io_x2; // @[MUL.scala 102:19]
  wire  m_1825_io_x3; // @[MUL.scala 102:19]
  wire  m_1825_io_s; // @[MUL.scala 102:19]
  wire  m_1825_io_cout; // @[MUL.scala 102:19]
  wire  m_1826_io_x1; // @[MUL.scala 102:19]
  wire  m_1826_io_x2; // @[MUL.scala 102:19]
  wire  m_1826_io_x3; // @[MUL.scala 102:19]
  wire  m_1826_io_s; // @[MUL.scala 102:19]
  wire  m_1826_io_cout; // @[MUL.scala 102:19]
  wire  m_1827_io_x1; // @[MUL.scala 102:19]
  wire  m_1827_io_x2; // @[MUL.scala 102:19]
  wire  m_1827_io_x3; // @[MUL.scala 102:19]
  wire  m_1827_io_s; // @[MUL.scala 102:19]
  wire  m_1827_io_cout; // @[MUL.scala 102:19]
  wire  m_1828_io_x1; // @[MUL.scala 102:19]
  wire  m_1828_io_x2; // @[MUL.scala 102:19]
  wire  m_1828_io_x3; // @[MUL.scala 102:19]
  wire  m_1828_io_s; // @[MUL.scala 102:19]
  wire  m_1828_io_cout; // @[MUL.scala 102:19]
  wire  m_1829_io_x1; // @[MUL.scala 102:19]
  wire  m_1829_io_x2; // @[MUL.scala 102:19]
  wire  m_1829_io_x3; // @[MUL.scala 102:19]
  wire  m_1829_io_s; // @[MUL.scala 102:19]
  wire  m_1829_io_cout; // @[MUL.scala 102:19]
  wire  m_1830_io_x1; // @[MUL.scala 102:19]
  wire  m_1830_io_x2; // @[MUL.scala 102:19]
  wire  m_1830_io_x3; // @[MUL.scala 102:19]
  wire  m_1830_io_s; // @[MUL.scala 102:19]
  wire  m_1830_io_cout; // @[MUL.scala 102:19]
  wire  m_1831_io_x1; // @[MUL.scala 102:19]
  wire  m_1831_io_x2; // @[MUL.scala 102:19]
  wire  m_1831_io_x3; // @[MUL.scala 102:19]
  wire  m_1831_io_s; // @[MUL.scala 102:19]
  wire  m_1831_io_cout; // @[MUL.scala 102:19]
  wire  m_1832_io_x1; // @[MUL.scala 102:19]
  wire  m_1832_io_x2; // @[MUL.scala 102:19]
  wire  m_1832_io_x3; // @[MUL.scala 102:19]
  wire  m_1832_io_s; // @[MUL.scala 102:19]
  wire  m_1832_io_cout; // @[MUL.scala 102:19]
  wire  m_1833_io_x1; // @[MUL.scala 102:19]
  wire  m_1833_io_x2; // @[MUL.scala 102:19]
  wire  m_1833_io_x3; // @[MUL.scala 102:19]
  wire  m_1833_io_s; // @[MUL.scala 102:19]
  wire  m_1833_io_cout; // @[MUL.scala 102:19]
  wire  m_1834_io_x1; // @[MUL.scala 102:19]
  wire  m_1834_io_x2; // @[MUL.scala 102:19]
  wire  m_1834_io_x3; // @[MUL.scala 102:19]
  wire  m_1834_io_s; // @[MUL.scala 102:19]
  wire  m_1834_io_cout; // @[MUL.scala 102:19]
  wire  m_1835_io_x1; // @[MUL.scala 102:19]
  wire  m_1835_io_x2; // @[MUL.scala 102:19]
  wire  m_1835_io_x3; // @[MUL.scala 102:19]
  wire  m_1835_io_s; // @[MUL.scala 102:19]
  wire  m_1835_io_cout; // @[MUL.scala 102:19]
  wire  m_1836_io_x1; // @[MUL.scala 102:19]
  wire  m_1836_io_x2; // @[MUL.scala 102:19]
  wire  m_1836_io_x3; // @[MUL.scala 102:19]
  wire  m_1836_io_s; // @[MUL.scala 102:19]
  wire  m_1836_io_cout; // @[MUL.scala 102:19]
  wire  m_1837_io_x1; // @[MUL.scala 102:19]
  wire  m_1837_io_x2; // @[MUL.scala 102:19]
  wire  m_1837_io_x3; // @[MUL.scala 102:19]
  wire  m_1837_io_s; // @[MUL.scala 102:19]
  wire  m_1837_io_cout; // @[MUL.scala 102:19]
  wire  m_1838_io_x1; // @[MUL.scala 102:19]
  wire  m_1838_io_x2; // @[MUL.scala 102:19]
  wire  m_1838_io_x3; // @[MUL.scala 102:19]
  wire  m_1838_io_s; // @[MUL.scala 102:19]
  wire  m_1838_io_cout; // @[MUL.scala 102:19]
  wire  m_1839_io_x1; // @[MUL.scala 102:19]
  wire  m_1839_io_x2; // @[MUL.scala 102:19]
  wire  m_1839_io_x3; // @[MUL.scala 102:19]
  wire  m_1839_io_s; // @[MUL.scala 102:19]
  wire  m_1839_io_cout; // @[MUL.scala 102:19]
  wire  m_1840_io_x1; // @[MUL.scala 102:19]
  wire  m_1840_io_x2; // @[MUL.scala 102:19]
  wire  m_1840_io_x3; // @[MUL.scala 102:19]
  wire  m_1840_io_s; // @[MUL.scala 102:19]
  wire  m_1840_io_cout; // @[MUL.scala 102:19]
  wire  m_1841_io_x1; // @[MUL.scala 102:19]
  wire  m_1841_io_x2; // @[MUL.scala 102:19]
  wire  m_1841_io_x3; // @[MUL.scala 102:19]
  wire  m_1841_io_s; // @[MUL.scala 102:19]
  wire  m_1841_io_cout; // @[MUL.scala 102:19]
  wire  m_1842_io_x1; // @[MUL.scala 102:19]
  wire  m_1842_io_x2; // @[MUL.scala 102:19]
  wire  m_1842_io_x3; // @[MUL.scala 102:19]
  wire  m_1842_io_s; // @[MUL.scala 102:19]
  wire  m_1842_io_cout; // @[MUL.scala 102:19]
  wire  m_1843_io_x1; // @[MUL.scala 102:19]
  wire  m_1843_io_x2; // @[MUL.scala 102:19]
  wire  m_1843_io_x3; // @[MUL.scala 102:19]
  wire  m_1843_io_s; // @[MUL.scala 102:19]
  wire  m_1843_io_cout; // @[MUL.scala 102:19]
  wire  m_1844_io_x1; // @[MUL.scala 102:19]
  wire  m_1844_io_x2; // @[MUL.scala 102:19]
  wire  m_1844_io_x3; // @[MUL.scala 102:19]
  wire  m_1844_io_s; // @[MUL.scala 102:19]
  wire  m_1844_io_cout; // @[MUL.scala 102:19]
  wire  m_1845_io_x1; // @[MUL.scala 102:19]
  wire  m_1845_io_x2; // @[MUL.scala 102:19]
  wire  m_1845_io_x3; // @[MUL.scala 102:19]
  wire  m_1845_io_s; // @[MUL.scala 102:19]
  wire  m_1845_io_cout; // @[MUL.scala 102:19]
  wire  m_1846_io_x1; // @[MUL.scala 102:19]
  wire  m_1846_io_x2; // @[MUL.scala 102:19]
  wire  m_1846_io_x3; // @[MUL.scala 102:19]
  wire  m_1846_io_s; // @[MUL.scala 102:19]
  wire  m_1846_io_cout; // @[MUL.scala 102:19]
  wire  m_1847_io_x1; // @[MUL.scala 102:19]
  wire  m_1847_io_x2; // @[MUL.scala 102:19]
  wire  m_1847_io_x3; // @[MUL.scala 102:19]
  wire  m_1847_io_s; // @[MUL.scala 102:19]
  wire  m_1847_io_cout; // @[MUL.scala 102:19]
  wire  m_1848_io_x1; // @[MUL.scala 102:19]
  wire  m_1848_io_x2; // @[MUL.scala 102:19]
  wire  m_1848_io_x3; // @[MUL.scala 102:19]
  wire  m_1848_io_s; // @[MUL.scala 102:19]
  wire  m_1848_io_cout; // @[MUL.scala 102:19]
  wire  m_1849_io_x1; // @[MUL.scala 102:19]
  wire  m_1849_io_x2; // @[MUL.scala 102:19]
  wire  m_1849_io_x3; // @[MUL.scala 102:19]
  wire  m_1849_io_s; // @[MUL.scala 102:19]
  wire  m_1849_io_cout; // @[MUL.scala 102:19]
  wire  m_1850_io_x1; // @[MUL.scala 102:19]
  wire  m_1850_io_x2; // @[MUL.scala 102:19]
  wire  m_1850_io_x3; // @[MUL.scala 102:19]
  wire  m_1850_io_s; // @[MUL.scala 102:19]
  wire  m_1850_io_cout; // @[MUL.scala 102:19]
  wire  m_1851_io_x1; // @[MUL.scala 102:19]
  wire  m_1851_io_x2; // @[MUL.scala 102:19]
  wire  m_1851_io_x3; // @[MUL.scala 102:19]
  wire  m_1851_io_s; // @[MUL.scala 102:19]
  wire  m_1851_io_cout; // @[MUL.scala 102:19]
  wire  m_1852_io_x1; // @[MUL.scala 102:19]
  wire  m_1852_io_x2; // @[MUL.scala 102:19]
  wire  m_1852_io_x3; // @[MUL.scala 102:19]
  wire  m_1852_io_s; // @[MUL.scala 102:19]
  wire  m_1852_io_cout; // @[MUL.scala 102:19]
  wire  m_1853_io_x1; // @[MUL.scala 102:19]
  wire  m_1853_io_x2; // @[MUL.scala 102:19]
  wire  m_1853_io_x3; // @[MUL.scala 102:19]
  wire  m_1853_io_s; // @[MUL.scala 102:19]
  wire  m_1853_io_cout; // @[MUL.scala 102:19]
  wire  m_1854_io_x1; // @[MUL.scala 102:19]
  wire  m_1854_io_x2; // @[MUL.scala 102:19]
  wire  m_1854_io_x3; // @[MUL.scala 102:19]
  wire  m_1854_io_s; // @[MUL.scala 102:19]
  wire  m_1854_io_cout; // @[MUL.scala 102:19]
  wire  m_1855_io_x1; // @[MUL.scala 102:19]
  wire  m_1855_io_x2; // @[MUL.scala 102:19]
  wire  m_1855_io_x3; // @[MUL.scala 102:19]
  wire  m_1855_io_s; // @[MUL.scala 102:19]
  wire  m_1855_io_cout; // @[MUL.scala 102:19]
  wire  m_1856_io_x1; // @[MUL.scala 102:19]
  wire  m_1856_io_x2; // @[MUL.scala 102:19]
  wire  m_1856_io_x3; // @[MUL.scala 102:19]
  wire  m_1856_io_s; // @[MUL.scala 102:19]
  wire  m_1856_io_cout; // @[MUL.scala 102:19]
  wire  m_1857_io_x1; // @[MUL.scala 102:19]
  wire  m_1857_io_x2; // @[MUL.scala 102:19]
  wire  m_1857_io_x3; // @[MUL.scala 102:19]
  wire  m_1857_io_s; // @[MUL.scala 102:19]
  wire  m_1857_io_cout; // @[MUL.scala 102:19]
  wire  m_1858_io_x1; // @[MUL.scala 102:19]
  wire  m_1858_io_x2; // @[MUL.scala 102:19]
  wire  m_1858_io_x3; // @[MUL.scala 102:19]
  wire  m_1858_io_s; // @[MUL.scala 102:19]
  wire  m_1858_io_cout; // @[MUL.scala 102:19]
  wire  m_1859_io_x1; // @[MUL.scala 102:19]
  wire  m_1859_io_x2; // @[MUL.scala 102:19]
  wire  m_1859_io_x3; // @[MUL.scala 102:19]
  wire  m_1859_io_s; // @[MUL.scala 102:19]
  wire  m_1859_io_cout; // @[MUL.scala 102:19]
  wire  m_1860_io_x1; // @[MUL.scala 102:19]
  wire  m_1860_io_x2; // @[MUL.scala 102:19]
  wire  m_1860_io_x3; // @[MUL.scala 102:19]
  wire  m_1860_io_s; // @[MUL.scala 102:19]
  wire  m_1860_io_cout; // @[MUL.scala 102:19]
  wire  m_1861_io_x1; // @[MUL.scala 102:19]
  wire  m_1861_io_x2; // @[MUL.scala 102:19]
  wire  m_1861_io_x3; // @[MUL.scala 102:19]
  wire  m_1861_io_s; // @[MUL.scala 102:19]
  wire  m_1861_io_cout; // @[MUL.scala 102:19]
  wire  m_1862_io_x1; // @[MUL.scala 102:19]
  wire  m_1862_io_x2; // @[MUL.scala 102:19]
  wire  m_1862_io_x3; // @[MUL.scala 102:19]
  wire  m_1862_io_s; // @[MUL.scala 102:19]
  wire  m_1862_io_cout; // @[MUL.scala 102:19]
  wire  m_1863_io_x1; // @[MUL.scala 102:19]
  wire  m_1863_io_x2; // @[MUL.scala 102:19]
  wire  m_1863_io_x3; // @[MUL.scala 102:19]
  wire  m_1863_io_s; // @[MUL.scala 102:19]
  wire  m_1863_io_cout; // @[MUL.scala 102:19]
  wire  m_1864_io_x1; // @[MUL.scala 102:19]
  wire  m_1864_io_x2; // @[MUL.scala 102:19]
  wire  m_1864_io_x3; // @[MUL.scala 102:19]
  wire  m_1864_io_s; // @[MUL.scala 102:19]
  wire  m_1864_io_cout; // @[MUL.scala 102:19]
  wire  m_1865_io_in_0; // @[MUL.scala 124:19]
  wire  m_1865_io_in_1; // @[MUL.scala 124:19]
  wire  m_1865_io_out_0; // @[MUL.scala 124:19]
  wire  m_1865_io_out_1; // @[MUL.scala 124:19]
  wire  m_1866_io_x1; // @[MUL.scala 102:19]
  wire  m_1866_io_x2; // @[MUL.scala 102:19]
  wire  m_1866_io_x3; // @[MUL.scala 102:19]
  wire  m_1866_io_s; // @[MUL.scala 102:19]
  wire  m_1866_io_cout; // @[MUL.scala 102:19]
  wire  m_1867_io_x1; // @[MUL.scala 102:19]
  wire  m_1867_io_x2; // @[MUL.scala 102:19]
  wire  m_1867_io_x3; // @[MUL.scala 102:19]
  wire  m_1867_io_s; // @[MUL.scala 102:19]
  wire  m_1867_io_cout; // @[MUL.scala 102:19]
  wire  m_1868_io_in_0; // @[MUL.scala 124:19]
  wire  m_1868_io_in_1; // @[MUL.scala 124:19]
  wire  m_1868_io_out_0; // @[MUL.scala 124:19]
  wire  m_1868_io_out_1; // @[MUL.scala 124:19]
  wire  m_1869_io_x1; // @[MUL.scala 102:19]
  wire  m_1869_io_x2; // @[MUL.scala 102:19]
  wire  m_1869_io_x3; // @[MUL.scala 102:19]
  wire  m_1869_io_s; // @[MUL.scala 102:19]
  wire  m_1869_io_cout; // @[MUL.scala 102:19]
  wire  m_1870_io_x1; // @[MUL.scala 102:19]
  wire  m_1870_io_x2; // @[MUL.scala 102:19]
  wire  m_1870_io_x3; // @[MUL.scala 102:19]
  wire  m_1870_io_s; // @[MUL.scala 102:19]
  wire  m_1870_io_cout; // @[MUL.scala 102:19]
  wire  m_1871_io_in_0; // @[MUL.scala 124:19]
  wire  m_1871_io_in_1; // @[MUL.scala 124:19]
  wire  m_1871_io_out_0; // @[MUL.scala 124:19]
  wire  m_1871_io_out_1; // @[MUL.scala 124:19]
  wire  m_1872_io_x1; // @[MUL.scala 102:19]
  wire  m_1872_io_x2; // @[MUL.scala 102:19]
  wire  m_1872_io_x3; // @[MUL.scala 102:19]
  wire  m_1872_io_s; // @[MUL.scala 102:19]
  wire  m_1872_io_cout; // @[MUL.scala 102:19]
  wire  m_1873_io_x1; // @[MUL.scala 102:19]
  wire  m_1873_io_x2; // @[MUL.scala 102:19]
  wire  m_1873_io_x3; // @[MUL.scala 102:19]
  wire  m_1873_io_s; // @[MUL.scala 102:19]
  wire  m_1873_io_cout; // @[MUL.scala 102:19]
  wire  m_1874_io_in_0; // @[MUL.scala 124:19]
  wire  m_1874_io_in_1; // @[MUL.scala 124:19]
  wire  m_1874_io_out_0; // @[MUL.scala 124:19]
  wire  m_1874_io_out_1; // @[MUL.scala 124:19]
  wire  m_1875_io_x1; // @[MUL.scala 102:19]
  wire  m_1875_io_x2; // @[MUL.scala 102:19]
  wire  m_1875_io_x3; // @[MUL.scala 102:19]
  wire  m_1875_io_s; // @[MUL.scala 102:19]
  wire  m_1875_io_cout; // @[MUL.scala 102:19]
  wire  m_1876_io_x1; // @[MUL.scala 102:19]
  wire  m_1876_io_x2; // @[MUL.scala 102:19]
  wire  m_1876_io_x3; // @[MUL.scala 102:19]
  wire  m_1876_io_s; // @[MUL.scala 102:19]
  wire  m_1876_io_cout; // @[MUL.scala 102:19]
  wire  m_1877_io_in_0; // @[MUL.scala 124:19]
  wire  m_1877_io_in_1; // @[MUL.scala 124:19]
  wire  m_1877_io_out_0; // @[MUL.scala 124:19]
  wire  m_1877_io_out_1; // @[MUL.scala 124:19]
  wire  m_1878_io_x1; // @[MUL.scala 102:19]
  wire  m_1878_io_x2; // @[MUL.scala 102:19]
  wire  m_1878_io_x3; // @[MUL.scala 102:19]
  wire  m_1878_io_s; // @[MUL.scala 102:19]
  wire  m_1878_io_cout; // @[MUL.scala 102:19]
  wire  m_1879_io_x1; // @[MUL.scala 102:19]
  wire  m_1879_io_x2; // @[MUL.scala 102:19]
  wire  m_1879_io_x3; // @[MUL.scala 102:19]
  wire  m_1879_io_s; // @[MUL.scala 102:19]
  wire  m_1879_io_cout; // @[MUL.scala 102:19]
  wire  m_1880_io_in_0; // @[MUL.scala 124:19]
  wire  m_1880_io_in_1; // @[MUL.scala 124:19]
  wire  m_1880_io_out_0; // @[MUL.scala 124:19]
  wire  m_1880_io_out_1; // @[MUL.scala 124:19]
  wire  m_1881_io_x1; // @[MUL.scala 102:19]
  wire  m_1881_io_x2; // @[MUL.scala 102:19]
  wire  m_1881_io_x3; // @[MUL.scala 102:19]
  wire  m_1881_io_s; // @[MUL.scala 102:19]
  wire  m_1881_io_cout; // @[MUL.scala 102:19]
  wire  m_1882_io_x1; // @[MUL.scala 102:19]
  wire  m_1882_io_x2; // @[MUL.scala 102:19]
  wire  m_1882_io_x3; // @[MUL.scala 102:19]
  wire  m_1882_io_s; // @[MUL.scala 102:19]
  wire  m_1882_io_cout; // @[MUL.scala 102:19]
  wire  m_1883_io_in_0; // @[MUL.scala 124:19]
  wire  m_1883_io_in_1; // @[MUL.scala 124:19]
  wire  m_1883_io_out_0; // @[MUL.scala 124:19]
  wire  m_1883_io_out_1; // @[MUL.scala 124:19]
  wire  m_1884_io_x1; // @[MUL.scala 102:19]
  wire  m_1884_io_x2; // @[MUL.scala 102:19]
  wire  m_1884_io_x3; // @[MUL.scala 102:19]
  wire  m_1884_io_s; // @[MUL.scala 102:19]
  wire  m_1884_io_cout; // @[MUL.scala 102:19]
  wire  m_1885_io_x1; // @[MUL.scala 102:19]
  wire  m_1885_io_x2; // @[MUL.scala 102:19]
  wire  m_1885_io_x3; // @[MUL.scala 102:19]
  wire  m_1885_io_s; // @[MUL.scala 102:19]
  wire  m_1885_io_cout; // @[MUL.scala 102:19]
  wire  m_1886_io_in_0; // @[MUL.scala 124:19]
  wire  m_1886_io_in_1; // @[MUL.scala 124:19]
  wire  m_1886_io_out_0; // @[MUL.scala 124:19]
  wire  m_1886_io_out_1; // @[MUL.scala 124:19]
  wire  m_1887_io_x1; // @[MUL.scala 102:19]
  wire  m_1887_io_x2; // @[MUL.scala 102:19]
  wire  m_1887_io_x3; // @[MUL.scala 102:19]
  wire  m_1887_io_s; // @[MUL.scala 102:19]
  wire  m_1887_io_cout; // @[MUL.scala 102:19]
  wire  m_1888_io_x1; // @[MUL.scala 102:19]
  wire  m_1888_io_x2; // @[MUL.scala 102:19]
  wire  m_1888_io_x3; // @[MUL.scala 102:19]
  wire  m_1888_io_s; // @[MUL.scala 102:19]
  wire  m_1888_io_cout; // @[MUL.scala 102:19]
  wire  m_1889_io_in_0; // @[MUL.scala 124:19]
  wire  m_1889_io_in_1; // @[MUL.scala 124:19]
  wire  m_1889_io_out_0; // @[MUL.scala 124:19]
  wire  m_1889_io_out_1; // @[MUL.scala 124:19]
  wire  m_1890_io_x1; // @[MUL.scala 102:19]
  wire  m_1890_io_x2; // @[MUL.scala 102:19]
  wire  m_1890_io_x3; // @[MUL.scala 102:19]
  wire  m_1890_io_s; // @[MUL.scala 102:19]
  wire  m_1890_io_cout; // @[MUL.scala 102:19]
  wire  m_1891_io_x1; // @[MUL.scala 102:19]
  wire  m_1891_io_x2; // @[MUL.scala 102:19]
  wire  m_1891_io_x3; // @[MUL.scala 102:19]
  wire  m_1891_io_s; // @[MUL.scala 102:19]
  wire  m_1891_io_cout; // @[MUL.scala 102:19]
  wire  m_1892_io_in_0; // @[MUL.scala 124:19]
  wire  m_1892_io_in_1; // @[MUL.scala 124:19]
  wire  m_1892_io_out_0; // @[MUL.scala 124:19]
  wire  m_1892_io_out_1; // @[MUL.scala 124:19]
  wire  m_1893_io_x1; // @[MUL.scala 102:19]
  wire  m_1893_io_x2; // @[MUL.scala 102:19]
  wire  m_1893_io_x3; // @[MUL.scala 102:19]
  wire  m_1893_io_s; // @[MUL.scala 102:19]
  wire  m_1893_io_cout; // @[MUL.scala 102:19]
  wire  m_1894_io_x1; // @[MUL.scala 102:19]
  wire  m_1894_io_x2; // @[MUL.scala 102:19]
  wire  m_1894_io_x3; // @[MUL.scala 102:19]
  wire  m_1894_io_s; // @[MUL.scala 102:19]
  wire  m_1894_io_cout; // @[MUL.scala 102:19]
  wire  m_1895_io_in_0; // @[MUL.scala 124:19]
  wire  m_1895_io_in_1; // @[MUL.scala 124:19]
  wire  m_1895_io_out_0; // @[MUL.scala 124:19]
  wire  m_1895_io_out_1; // @[MUL.scala 124:19]
  wire  m_1896_io_x1; // @[MUL.scala 102:19]
  wire  m_1896_io_x2; // @[MUL.scala 102:19]
  wire  m_1896_io_x3; // @[MUL.scala 102:19]
  wire  m_1896_io_s; // @[MUL.scala 102:19]
  wire  m_1896_io_cout; // @[MUL.scala 102:19]
  wire  m_1897_io_x1; // @[MUL.scala 102:19]
  wire  m_1897_io_x2; // @[MUL.scala 102:19]
  wire  m_1897_io_x3; // @[MUL.scala 102:19]
  wire  m_1897_io_s; // @[MUL.scala 102:19]
  wire  m_1897_io_cout; // @[MUL.scala 102:19]
  wire  m_1898_io_x1; // @[MUL.scala 102:19]
  wire  m_1898_io_x2; // @[MUL.scala 102:19]
  wire  m_1898_io_x3; // @[MUL.scala 102:19]
  wire  m_1898_io_s; // @[MUL.scala 102:19]
  wire  m_1898_io_cout; // @[MUL.scala 102:19]
  wire  m_1899_io_x1; // @[MUL.scala 102:19]
  wire  m_1899_io_x2; // @[MUL.scala 102:19]
  wire  m_1899_io_x3; // @[MUL.scala 102:19]
  wire  m_1899_io_s; // @[MUL.scala 102:19]
  wire  m_1899_io_cout; // @[MUL.scala 102:19]
  wire  m_1900_io_x1; // @[MUL.scala 102:19]
  wire  m_1900_io_x2; // @[MUL.scala 102:19]
  wire  m_1900_io_x3; // @[MUL.scala 102:19]
  wire  m_1900_io_s; // @[MUL.scala 102:19]
  wire  m_1900_io_cout; // @[MUL.scala 102:19]
  wire  m_1901_io_x1; // @[MUL.scala 102:19]
  wire  m_1901_io_x2; // @[MUL.scala 102:19]
  wire  m_1901_io_x3; // @[MUL.scala 102:19]
  wire  m_1901_io_s; // @[MUL.scala 102:19]
  wire  m_1901_io_cout; // @[MUL.scala 102:19]
  wire  m_1902_io_x1; // @[MUL.scala 102:19]
  wire  m_1902_io_x2; // @[MUL.scala 102:19]
  wire  m_1902_io_x3; // @[MUL.scala 102:19]
  wire  m_1902_io_s; // @[MUL.scala 102:19]
  wire  m_1902_io_cout; // @[MUL.scala 102:19]
  wire  m_1903_io_x1; // @[MUL.scala 102:19]
  wire  m_1903_io_x2; // @[MUL.scala 102:19]
  wire  m_1903_io_x3; // @[MUL.scala 102:19]
  wire  m_1903_io_s; // @[MUL.scala 102:19]
  wire  m_1903_io_cout; // @[MUL.scala 102:19]
  wire  m_1904_io_x1; // @[MUL.scala 102:19]
  wire  m_1904_io_x2; // @[MUL.scala 102:19]
  wire  m_1904_io_x3; // @[MUL.scala 102:19]
  wire  m_1904_io_s; // @[MUL.scala 102:19]
  wire  m_1904_io_cout; // @[MUL.scala 102:19]
  wire  m_1905_io_x1; // @[MUL.scala 102:19]
  wire  m_1905_io_x2; // @[MUL.scala 102:19]
  wire  m_1905_io_x3; // @[MUL.scala 102:19]
  wire  m_1905_io_s; // @[MUL.scala 102:19]
  wire  m_1905_io_cout; // @[MUL.scala 102:19]
  wire  m_1906_io_x1; // @[MUL.scala 102:19]
  wire  m_1906_io_x2; // @[MUL.scala 102:19]
  wire  m_1906_io_x3; // @[MUL.scala 102:19]
  wire  m_1906_io_s; // @[MUL.scala 102:19]
  wire  m_1906_io_cout; // @[MUL.scala 102:19]
  wire  m_1907_io_x1; // @[MUL.scala 102:19]
  wire  m_1907_io_x2; // @[MUL.scala 102:19]
  wire  m_1907_io_x3; // @[MUL.scala 102:19]
  wire  m_1907_io_s; // @[MUL.scala 102:19]
  wire  m_1907_io_cout; // @[MUL.scala 102:19]
  wire  m_1908_io_x1; // @[MUL.scala 102:19]
  wire  m_1908_io_x2; // @[MUL.scala 102:19]
  wire  m_1908_io_x3; // @[MUL.scala 102:19]
  wire  m_1908_io_s; // @[MUL.scala 102:19]
  wire  m_1908_io_cout; // @[MUL.scala 102:19]
  wire  m_1909_io_x1; // @[MUL.scala 102:19]
  wire  m_1909_io_x2; // @[MUL.scala 102:19]
  wire  m_1909_io_x3; // @[MUL.scala 102:19]
  wire  m_1909_io_s; // @[MUL.scala 102:19]
  wire  m_1909_io_cout; // @[MUL.scala 102:19]
  wire  m_1910_io_x1; // @[MUL.scala 102:19]
  wire  m_1910_io_x2; // @[MUL.scala 102:19]
  wire  m_1910_io_x3; // @[MUL.scala 102:19]
  wire  m_1910_io_s; // @[MUL.scala 102:19]
  wire  m_1910_io_cout; // @[MUL.scala 102:19]
  wire  m_1911_io_x1; // @[MUL.scala 102:19]
  wire  m_1911_io_x2; // @[MUL.scala 102:19]
  wire  m_1911_io_x3; // @[MUL.scala 102:19]
  wire  m_1911_io_s; // @[MUL.scala 102:19]
  wire  m_1911_io_cout; // @[MUL.scala 102:19]
  wire  m_1912_io_x1; // @[MUL.scala 102:19]
  wire  m_1912_io_x2; // @[MUL.scala 102:19]
  wire  m_1912_io_x3; // @[MUL.scala 102:19]
  wire  m_1912_io_s; // @[MUL.scala 102:19]
  wire  m_1912_io_cout; // @[MUL.scala 102:19]
  wire  m_1913_io_x1; // @[MUL.scala 102:19]
  wire  m_1913_io_x2; // @[MUL.scala 102:19]
  wire  m_1913_io_x3; // @[MUL.scala 102:19]
  wire  m_1913_io_s; // @[MUL.scala 102:19]
  wire  m_1913_io_cout; // @[MUL.scala 102:19]
  wire  m_1914_io_x1; // @[MUL.scala 102:19]
  wire  m_1914_io_x2; // @[MUL.scala 102:19]
  wire  m_1914_io_x3; // @[MUL.scala 102:19]
  wire  m_1914_io_s; // @[MUL.scala 102:19]
  wire  m_1914_io_cout; // @[MUL.scala 102:19]
  wire  m_1915_io_x1; // @[MUL.scala 102:19]
  wire  m_1915_io_x2; // @[MUL.scala 102:19]
  wire  m_1915_io_x3; // @[MUL.scala 102:19]
  wire  m_1915_io_s; // @[MUL.scala 102:19]
  wire  m_1915_io_cout; // @[MUL.scala 102:19]
  wire  m_1916_io_x1; // @[MUL.scala 102:19]
  wire  m_1916_io_x2; // @[MUL.scala 102:19]
  wire  m_1916_io_x3; // @[MUL.scala 102:19]
  wire  m_1916_io_s; // @[MUL.scala 102:19]
  wire  m_1916_io_cout; // @[MUL.scala 102:19]
  wire  m_1917_io_x1; // @[MUL.scala 102:19]
  wire  m_1917_io_x2; // @[MUL.scala 102:19]
  wire  m_1917_io_x3; // @[MUL.scala 102:19]
  wire  m_1917_io_s; // @[MUL.scala 102:19]
  wire  m_1917_io_cout; // @[MUL.scala 102:19]
  wire  m_1918_io_x1; // @[MUL.scala 102:19]
  wire  m_1918_io_x2; // @[MUL.scala 102:19]
  wire  m_1918_io_x3; // @[MUL.scala 102:19]
  wire  m_1918_io_s; // @[MUL.scala 102:19]
  wire  m_1918_io_cout; // @[MUL.scala 102:19]
  wire  m_1919_io_x1; // @[MUL.scala 102:19]
  wire  m_1919_io_x2; // @[MUL.scala 102:19]
  wire  m_1919_io_x3; // @[MUL.scala 102:19]
  wire  m_1919_io_s; // @[MUL.scala 102:19]
  wire  m_1919_io_cout; // @[MUL.scala 102:19]
  wire  m_1920_io_x1; // @[MUL.scala 102:19]
  wire  m_1920_io_x2; // @[MUL.scala 102:19]
  wire  m_1920_io_x3; // @[MUL.scala 102:19]
  wire  m_1920_io_s; // @[MUL.scala 102:19]
  wire  m_1920_io_cout; // @[MUL.scala 102:19]
  wire  m_1921_io_x1; // @[MUL.scala 102:19]
  wire  m_1921_io_x2; // @[MUL.scala 102:19]
  wire  m_1921_io_x3; // @[MUL.scala 102:19]
  wire  m_1921_io_s; // @[MUL.scala 102:19]
  wire  m_1921_io_cout; // @[MUL.scala 102:19]
  wire  m_1922_io_x1; // @[MUL.scala 102:19]
  wire  m_1922_io_x2; // @[MUL.scala 102:19]
  wire  m_1922_io_x3; // @[MUL.scala 102:19]
  wire  m_1922_io_s; // @[MUL.scala 102:19]
  wire  m_1922_io_cout; // @[MUL.scala 102:19]
  wire  m_1923_io_x1; // @[MUL.scala 102:19]
  wire  m_1923_io_x2; // @[MUL.scala 102:19]
  wire  m_1923_io_x3; // @[MUL.scala 102:19]
  wire  m_1923_io_s; // @[MUL.scala 102:19]
  wire  m_1923_io_cout; // @[MUL.scala 102:19]
  wire  m_1924_io_x1; // @[MUL.scala 102:19]
  wire  m_1924_io_x2; // @[MUL.scala 102:19]
  wire  m_1924_io_x3; // @[MUL.scala 102:19]
  wire  m_1924_io_s; // @[MUL.scala 102:19]
  wire  m_1924_io_cout; // @[MUL.scala 102:19]
  wire  m_1925_io_in_0; // @[MUL.scala 124:19]
  wire  m_1925_io_in_1; // @[MUL.scala 124:19]
  wire  m_1925_io_out_0; // @[MUL.scala 124:19]
  wire  m_1925_io_out_1; // @[MUL.scala 124:19]
  wire  m_1926_io_x1; // @[MUL.scala 102:19]
  wire  m_1926_io_x2; // @[MUL.scala 102:19]
  wire  m_1926_io_x3; // @[MUL.scala 102:19]
  wire  m_1926_io_s; // @[MUL.scala 102:19]
  wire  m_1926_io_cout; // @[MUL.scala 102:19]
  wire  m_1927_io_in_0; // @[MUL.scala 124:19]
  wire  m_1927_io_in_1; // @[MUL.scala 124:19]
  wire  m_1927_io_out_0; // @[MUL.scala 124:19]
  wire  m_1927_io_out_1; // @[MUL.scala 124:19]
  wire  m_1928_io_x1; // @[MUL.scala 102:19]
  wire  m_1928_io_x2; // @[MUL.scala 102:19]
  wire  m_1928_io_x3; // @[MUL.scala 102:19]
  wire  m_1928_io_s; // @[MUL.scala 102:19]
  wire  m_1928_io_cout; // @[MUL.scala 102:19]
  wire  m_1929_io_in_0; // @[MUL.scala 124:19]
  wire  m_1929_io_in_1; // @[MUL.scala 124:19]
  wire  m_1929_io_out_0; // @[MUL.scala 124:19]
  wire  m_1929_io_out_1; // @[MUL.scala 124:19]
  wire  m_1930_io_x1; // @[MUL.scala 102:19]
  wire  m_1930_io_x2; // @[MUL.scala 102:19]
  wire  m_1930_io_x3; // @[MUL.scala 102:19]
  wire  m_1930_io_s; // @[MUL.scala 102:19]
  wire  m_1930_io_cout; // @[MUL.scala 102:19]
  wire  m_1931_io_x1; // @[MUL.scala 102:19]
  wire  m_1931_io_x2; // @[MUL.scala 102:19]
  wire  m_1931_io_x3; // @[MUL.scala 102:19]
  wire  m_1931_io_s; // @[MUL.scala 102:19]
  wire  m_1931_io_cout; // @[MUL.scala 102:19]
  wire  m_1932_io_x1; // @[MUL.scala 102:19]
  wire  m_1932_io_x2; // @[MUL.scala 102:19]
  wire  m_1932_io_x3; // @[MUL.scala 102:19]
  wire  m_1932_io_s; // @[MUL.scala 102:19]
  wire  m_1932_io_cout; // @[MUL.scala 102:19]
  wire  m_1933_io_x1; // @[MUL.scala 102:19]
  wire  m_1933_io_x2; // @[MUL.scala 102:19]
  wire  m_1933_io_x3; // @[MUL.scala 102:19]
  wire  m_1933_io_s; // @[MUL.scala 102:19]
  wire  m_1933_io_cout; // @[MUL.scala 102:19]
  wire  m_1934_io_x1; // @[MUL.scala 102:19]
  wire  m_1934_io_x2; // @[MUL.scala 102:19]
  wire  m_1934_io_x3; // @[MUL.scala 102:19]
  wire  m_1934_io_s; // @[MUL.scala 102:19]
  wire  m_1934_io_cout; // @[MUL.scala 102:19]
  wire  m_1935_io_x1; // @[MUL.scala 102:19]
  wire  m_1935_io_x2; // @[MUL.scala 102:19]
  wire  m_1935_io_x3; // @[MUL.scala 102:19]
  wire  m_1935_io_s; // @[MUL.scala 102:19]
  wire  m_1935_io_cout; // @[MUL.scala 102:19]
  wire  m_1936_io_x1; // @[MUL.scala 102:19]
  wire  m_1936_io_x2; // @[MUL.scala 102:19]
  wire  m_1936_io_x3; // @[MUL.scala 102:19]
  wire  m_1936_io_s; // @[MUL.scala 102:19]
  wire  m_1936_io_cout; // @[MUL.scala 102:19]
  wire  m_1937_io_x1; // @[MUL.scala 102:19]
  wire  m_1937_io_x2; // @[MUL.scala 102:19]
  wire  m_1937_io_x3; // @[MUL.scala 102:19]
  wire  m_1937_io_s; // @[MUL.scala 102:19]
  wire  m_1937_io_cout; // @[MUL.scala 102:19]
  wire  m_1938_io_x1; // @[MUL.scala 102:19]
  wire  m_1938_io_x2; // @[MUL.scala 102:19]
  wire  m_1938_io_x3; // @[MUL.scala 102:19]
  wire  m_1938_io_s; // @[MUL.scala 102:19]
  wire  m_1938_io_cout; // @[MUL.scala 102:19]
  wire  m_1939_io_x1; // @[MUL.scala 102:19]
  wire  m_1939_io_x2; // @[MUL.scala 102:19]
  wire  m_1939_io_x3; // @[MUL.scala 102:19]
  wire  m_1939_io_s; // @[MUL.scala 102:19]
  wire  m_1939_io_cout; // @[MUL.scala 102:19]
  wire  m_1940_io_x1; // @[MUL.scala 102:19]
  wire  m_1940_io_x2; // @[MUL.scala 102:19]
  wire  m_1940_io_x3; // @[MUL.scala 102:19]
  wire  m_1940_io_s; // @[MUL.scala 102:19]
  wire  m_1940_io_cout; // @[MUL.scala 102:19]
  wire  m_1941_io_x1; // @[MUL.scala 102:19]
  wire  m_1941_io_x2; // @[MUL.scala 102:19]
  wire  m_1941_io_x3; // @[MUL.scala 102:19]
  wire  m_1941_io_s; // @[MUL.scala 102:19]
  wire  m_1941_io_cout; // @[MUL.scala 102:19]
  wire  m_1942_io_x1; // @[MUL.scala 102:19]
  wire  m_1942_io_x2; // @[MUL.scala 102:19]
  wire  m_1942_io_x3; // @[MUL.scala 102:19]
  wire  m_1942_io_s; // @[MUL.scala 102:19]
  wire  m_1942_io_cout; // @[MUL.scala 102:19]
  wire  m_1943_io_x1; // @[MUL.scala 102:19]
  wire  m_1943_io_x2; // @[MUL.scala 102:19]
  wire  m_1943_io_x3; // @[MUL.scala 102:19]
  wire  m_1943_io_s; // @[MUL.scala 102:19]
  wire  m_1943_io_cout; // @[MUL.scala 102:19]
  wire  m_1944_io_in_0; // @[MUL.scala 124:19]
  wire  m_1944_io_in_1; // @[MUL.scala 124:19]
  wire  m_1944_io_out_0; // @[MUL.scala 124:19]
  wire  m_1944_io_out_1; // @[MUL.scala 124:19]
  wire  m_1945_io_in_0; // @[MUL.scala 124:19]
  wire  m_1945_io_in_1; // @[MUL.scala 124:19]
  wire  m_1945_io_out_0; // @[MUL.scala 124:19]
  wire  m_1945_io_out_1; // @[MUL.scala 124:19]
  wire  m_1946_io_in_0; // @[MUL.scala 124:19]
  wire  m_1946_io_in_1; // @[MUL.scala 124:19]
  wire  m_1946_io_out_0; // @[MUL.scala 124:19]
  wire  m_1946_io_out_1; // @[MUL.scala 124:19]
  wire  m_1947_io_in_0; // @[MUL.scala 124:19]
  wire  m_1947_io_in_1; // @[MUL.scala 124:19]
  wire  m_1947_io_out_0; // @[MUL.scala 124:19]
  wire  m_1947_io_out_1; // @[MUL.scala 124:19]
  wire  m_1948_io_in_0; // @[MUL.scala 124:19]
  wire  m_1948_io_in_1; // @[MUL.scala 124:19]
  wire  m_1948_io_out_0; // @[MUL.scala 124:19]
  wire  m_1948_io_out_1; // @[MUL.scala 124:19]
  wire  m_1949_io_in_0; // @[MUL.scala 124:19]
  wire  m_1949_io_in_1; // @[MUL.scala 124:19]
  wire  m_1949_io_out_0; // @[MUL.scala 124:19]
  wire  m_1949_io_out_1; // @[MUL.scala 124:19]
  wire  m_1950_io_in_0; // @[MUL.scala 124:19]
  wire  m_1950_io_in_1; // @[MUL.scala 124:19]
  wire  m_1950_io_out_0; // @[MUL.scala 124:19]
  wire  m_1950_io_out_1; // @[MUL.scala 124:19]
  wire  m_1951_io_in_0; // @[MUL.scala 124:19]
  wire  m_1951_io_in_1; // @[MUL.scala 124:19]
  wire  m_1951_io_out_0; // @[MUL.scala 124:19]
  wire  m_1951_io_out_1; // @[MUL.scala 124:19]
  wire  m_1952_io_in_0; // @[MUL.scala 124:19]
  wire  m_1952_io_in_1; // @[MUL.scala 124:19]
  wire  m_1952_io_out_0; // @[MUL.scala 124:19]
  wire  m_1952_io_out_1; // @[MUL.scala 124:19]
  wire  m_1953_io_in_0; // @[MUL.scala 124:19]
  wire  m_1953_io_in_1; // @[MUL.scala 124:19]
  wire  m_1953_io_out_0; // @[MUL.scala 124:19]
  wire  m_1953_io_out_1; // @[MUL.scala 124:19]
  wire  m_1954_io_in_0; // @[MUL.scala 124:19]
  wire  m_1954_io_in_1; // @[MUL.scala 124:19]
  wire  m_1954_io_out_0; // @[MUL.scala 124:19]
  wire  m_1954_io_out_1; // @[MUL.scala 124:19]
  wire  m_1955_io_in_0; // @[MUL.scala 124:19]
  wire  m_1955_io_in_1; // @[MUL.scala 124:19]
  wire  m_1955_io_out_0; // @[MUL.scala 124:19]
  wire  m_1955_io_out_1; // @[MUL.scala 124:19]
  wire  m_1956_io_in_0; // @[MUL.scala 124:19]
  wire  m_1956_io_in_1; // @[MUL.scala 124:19]
  wire  m_1956_io_out_0; // @[MUL.scala 124:19]
  wire  m_1956_io_out_1; // @[MUL.scala 124:19]
  wire  m_1957_io_in_0; // @[MUL.scala 124:19]
  wire  m_1957_io_in_1; // @[MUL.scala 124:19]
  wire  m_1957_io_out_0; // @[MUL.scala 124:19]
  wire  m_1957_io_out_1; // @[MUL.scala 124:19]
  wire  m_1958_io_in_0; // @[MUL.scala 124:19]
  wire  m_1958_io_in_1; // @[MUL.scala 124:19]
  wire  m_1958_io_out_0; // @[MUL.scala 124:19]
  wire  m_1958_io_out_1; // @[MUL.scala 124:19]
  wire  m_1959_io_in_0; // @[MUL.scala 124:19]
  wire  m_1959_io_in_1; // @[MUL.scala 124:19]
  wire  m_1959_io_out_0; // @[MUL.scala 124:19]
  wire  m_1959_io_out_1; // @[MUL.scala 124:19]
  wire  m_1960_io_in_0; // @[MUL.scala 124:19]
  wire  m_1960_io_in_1; // @[MUL.scala 124:19]
  wire  m_1960_io_out_0; // @[MUL.scala 124:19]
  wire  m_1960_io_out_1; // @[MUL.scala 124:19]
  wire  m_1961_io_in_0; // @[MUL.scala 124:19]
  wire  m_1961_io_in_1; // @[MUL.scala 124:19]
  wire  m_1961_io_out_0; // @[MUL.scala 124:19]
  wire  m_1961_io_out_1; // @[MUL.scala 124:19]
  wire  m_1962_io_in_0; // @[MUL.scala 124:19]
  wire  m_1962_io_in_1; // @[MUL.scala 124:19]
  wire  m_1962_io_out_0; // @[MUL.scala 124:19]
  wire  m_1962_io_out_1; // @[MUL.scala 124:19]
  wire  m_1963_io_in_0; // @[MUL.scala 124:19]
  wire  m_1963_io_in_1; // @[MUL.scala 124:19]
  wire  m_1963_io_out_0; // @[MUL.scala 124:19]
  wire  m_1963_io_out_1; // @[MUL.scala 124:19]
  wire  m_1964_io_in_0; // @[MUL.scala 124:19]
  wire  m_1964_io_in_1; // @[MUL.scala 124:19]
  wire  m_1964_io_out_0; // @[MUL.scala 124:19]
  wire  m_1964_io_out_1; // @[MUL.scala 124:19]
  wire  m_1965_io_in_0; // @[MUL.scala 124:19]
  wire  m_1965_io_in_1; // @[MUL.scala 124:19]
  wire  m_1965_io_out_0; // @[MUL.scala 124:19]
  wire  m_1965_io_out_1; // @[MUL.scala 124:19]
  wire  m_1966_io_in_0; // @[MUL.scala 124:19]
  wire  m_1966_io_in_1; // @[MUL.scala 124:19]
  wire  m_1966_io_out_0; // @[MUL.scala 124:19]
  wire  m_1966_io_out_1; // @[MUL.scala 124:19]
  wire  m_1967_io_x1; // @[MUL.scala 102:19]
  wire  m_1967_io_x2; // @[MUL.scala 102:19]
  wire  m_1967_io_x3; // @[MUL.scala 102:19]
  wire  m_1967_io_s; // @[MUL.scala 102:19]
  wire  m_1967_io_cout; // @[MUL.scala 102:19]
  wire  m_1968_io_x1; // @[MUL.scala 102:19]
  wire  m_1968_io_x2; // @[MUL.scala 102:19]
  wire  m_1968_io_x3; // @[MUL.scala 102:19]
  wire  m_1968_io_s; // @[MUL.scala 102:19]
  wire  m_1968_io_cout; // @[MUL.scala 102:19]
  wire  m_1969_io_x1; // @[MUL.scala 102:19]
  wire  m_1969_io_x2; // @[MUL.scala 102:19]
  wire  m_1969_io_x3; // @[MUL.scala 102:19]
  wire  m_1969_io_s; // @[MUL.scala 102:19]
  wire  m_1969_io_cout; // @[MUL.scala 102:19]
  wire  m_1970_io_x1; // @[MUL.scala 102:19]
  wire  m_1970_io_x2; // @[MUL.scala 102:19]
  wire  m_1970_io_x3; // @[MUL.scala 102:19]
  wire  m_1970_io_s; // @[MUL.scala 102:19]
  wire  m_1970_io_cout; // @[MUL.scala 102:19]
  wire  m_1971_io_x1; // @[MUL.scala 102:19]
  wire  m_1971_io_x2; // @[MUL.scala 102:19]
  wire  m_1971_io_x3; // @[MUL.scala 102:19]
  wire  m_1971_io_s; // @[MUL.scala 102:19]
  wire  m_1971_io_cout; // @[MUL.scala 102:19]
  wire  m_1972_io_x1; // @[MUL.scala 102:19]
  wire  m_1972_io_x2; // @[MUL.scala 102:19]
  wire  m_1972_io_x3; // @[MUL.scala 102:19]
  wire  m_1972_io_s; // @[MUL.scala 102:19]
  wire  m_1972_io_cout; // @[MUL.scala 102:19]
  wire  m_1973_io_x1; // @[MUL.scala 102:19]
  wire  m_1973_io_x2; // @[MUL.scala 102:19]
  wire  m_1973_io_x3; // @[MUL.scala 102:19]
  wire  m_1973_io_s; // @[MUL.scala 102:19]
  wire  m_1973_io_cout; // @[MUL.scala 102:19]
  wire  m_1974_io_x1; // @[MUL.scala 102:19]
  wire  m_1974_io_x2; // @[MUL.scala 102:19]
  wire  m_1974_io_x3; // @[MUL.scala 102:19]
  wire  m_1974_io_s; // @[MUL.scala 102:19]
  wire  m_1974_io_cout; // @[MUL.scala 102:19]
  wire  m_1975_io_x1; // @[MUL.scala 102:19]
  wire  m_1975_io_x2; // @[MUL.scala 102:19]
  wire  m_1975_io_x3; // @[MUL.scala 102:19]
  wire  m_1975_io_s; // @[MUL.scala 102:19]
  wire  m_1975_io_cout; // @[MUL.scala 102:19]
  wire  m_1976_io_x1; // @[MUL.scala 102:19]
  wire  m_1976_io_x2; // @[MUL.scala 102:19]
  wire  m_1976_io_x3; // @[MUL.scala 102:19]
  wire  m_1976_io_s; // @[MUL.scala 102:19]
  wire  m_1976_io_cout; // @[MUL.scala 102:19]
  wire  m_1977_io_x1; // @[MUL.scala 102:19]
  wire  m_1977_io_x2; // @[MUL.scala 102:19]
  wire  m_1977_io_x3; // @[MUL.scala 102:19]
  wire  m_1977_io_s; // @[MUL.scala 102:19]
  wire  m_1977_io_cout; // @[MUL.scala 102:19]
  wire  m_1978_io_x1; // @[MUL.scala 102:19]
  wire  m_1978_io_x2; // @[MUL.scala 102:19]
  wire  m_1978_io_x3; // @[MUL.scala 102:19]
  wire  m_1978_io_s; // @[MUL.scala 102:19]
  wire  m_1978_io_cout; // @[MUL.scala 102:19]
  wire  m_1979_io_x1; // @[MUL.scala 102:19]
  wire  m_1979_io_x2; // @[MUL.scala 102:19]
  wire  m_1979_io_x3; // @[MUL.scala 102:19]
  wire  m_1979_io_s; // @[MUL.scala 102:19]
  wire  m_1979_io_cout; // @[MUL.scala 102:19]
  wire  m_1980_io_x1; // @[MUL.scala 102:19]
  wire  m_1980_io_x2; // @[MUL.scala 102:19]
  wire  m_1980_io_x3; // @[MUL.scala 102:19]
  wire  m_1980_io_s; // @[MUL.scala 102:19]
  wire  m_1980_io_cout; // @[MUL.scala 102:19]
  wire  m_1981_io_x1; // @[MUL.scala 102:19]
  wire  m_1981_io_x2; // @[MUL.scala 102:19]
  wire  m_1981_io_x3; // @[MUL.scala 102:19]
  wire  m_1981_io_s; // @[MUL.scala 102:19]
  wire  m_1981_io_cout; // @[MUL.scala 102:19]
  wire  m_1982_io_x1; // @[MUL.scala 102:19]
  wire  m_1982_io_x2; // @[MUL.scala 102:19]
  wire  m_1982_io_x3; // @[MUL.scala 102:19]
  wire  m_1982_io_s; // @[MUL.scala 102:19]
  wire  m_1982_io_cout; // @[MUL.scala 102:19]
  wire  m_1983_io_x1; // @[MUL.scala 102:19]
  wire  m_1983_io_x2; // @[MUL.scala 102:19]
  wire  m_1983_io_x3; // @[MUL.scala 102:19]
  wire  m_1983_io_s; // @[MUL.scala 102:19]
  wire  m_1983_io_cout; // @[MUL.scala 102:19]
  wire  m_1984_io_x1; // @[MUL.scala 102:19]
  wire  m_1984_io_x2; // @[MUL.scala 102:19]
  wire  m_1984_io_x3; // @[MUL.scala 102:19]
  wire  m_1984_io_s; // @[MUL.scala 102:19]
  wire  m_1984_io_cout; // @[MUL.scala 102:19]
  wire  m_1985_io_x1; // @[MUL.scala 102:19]
  wire  m_1985_io_x2; // @[MUL.scala 102:19]
  wire  m_1985_io_x3; // @[MUL.scala 102:19]
  wire  m_1985_io_s; // @[MUL.scala 102:19]
  wire  m_1985_io_cout; // @[MUL.scala 102:19]
  wire  m_1986_io_x1; // @[MUL.scala 102:19]
  wire  m_1986_io_x2; // @[MUL.scala 102:19]
  wire  m_1986_io_x3; // @[MUL.scala 102:19]
  wire  m_1986_io_s; // @[MUL.scala 102:19]
  wire  m_1986_io_cout; // @[MUL.scala 102:19]
  wire  m_1987_io_x1; // @[MUL.scala 102:19]
  wire  m_1987_io_x2; // @[MUL.scala 102:19]
  wire  m_1987_io_x3; // @[MUL.scala 102:19]
  wire  m_1987_io_s; // @[MUL.scala 102:19]
  wire  m_1987_io_cout; // @[MUL.scala 102:19]
  wire  m_1988_io_x1; // @[MUL.scala 102:19]
  wire  m_1988_io_x2; // @[MUL.scala 102:19]
  wire  m_1988_io_x3; // @[MUL.scala 102:19]
  wire  m_1988_io_s; // @[MUL.scala 102:19]
  wire  m_1988_io_cout; // @[MUL.scala 102:19]
  wire  m_1989_io_in_0; // @[MUL.scala 124:19]
  wire  m_1989_io_in_1; // @[MUL.scala 124:19]
  wire  m_1989_io_out_0; // @[MUL.scala 124:19]
  wire  m_1989_io_out_1; // @[MUL.scala 124:19]
  wire  m_1990_io_x1; // @[MUL.scala 102:19]
  wire  m_1990_io_x2; // @[MUL.scala 102:19]
  wire  m_1990_io_x3; // @[MUL.scala 102:19]
  wire  m_1990_io_s; // @[MUL.scala 102:19]
  wire  m_1990_io_cout; // @[MUL.scala 102:19]
  wire  m_1991_io_in_0; // @[MUL.scala 124:19]
  wire  m_1991_io_in_1; // @[MUL.scala 124:19]
  wire  m_1991_io_out_0; // @[MUL.scala 124:19]
  wire  m_1991_io_out_1; // @[MUL.scala 124:19]
  wire  m_1992_io_x1; // @[MUL.scala 102:19]
  wire  m_1992_io_x2; // @[MUL.scala 102:19]
  wire  m_1992_io_x3; // @[MUL.scala 102:19]
  wire  m_1992_io_s; // @[MUL.scala 102:19]
  wire  m_1992_io_cout; // @[MUL.scala 102:19]
  wire  m_1993_io_in_0; // @[MUL.scala 124:19]
  wire  m_1993_io_in_1; // @[MUL.scala 124:19]
  wire  m_1993_io_out_0; // @[MUL.scala 124:19]
  wire  m_1993_io_out_1; // @[MUL.scala 124:19]
  wire  m_1994_io_x1; // @[MUL.scala 102:19]
  wire  m_1994_io_x2; // @[MUL.scala 102:19]
  wire  m_1994_io_x3; // @[MUL.scala 102:19]
  wire  m_1994_io_s; // @[MUL.scala 102:19]
  wire  m_1994_io_cout; // @[MUL.scala 102:19]
  wire  m_1995_io_in_0; // @[MUL.scala 124:19]
  wire  m_1995_io_in_1; // @[MUL.scala 124:19]
  wire  m_1995_io_out_0; // @[MUL.scala 124:19]
  wire  m_1995_io_out_1; // @[MUL.scala 124:19]
  wire  m_1996_io_x1; // @[MUL.scala 102:19]
  wire  m_1996_io_x2; // @[MUL.scala 102:19]
  wire  m_1996_io_x3; // @[MUL.scala 102:19]
  wire  m_1996_io_s; // @[MUL.scala 102:19]
  wire  m_1996_io_cout; // @[MUL.scala 102:19]
  wire  m_1997_io_in_0; // @[MUL.scala 124:19]
  wire  m_1997_io_in_1; // @[MUL.scala 124:19]
  wire  m_1997_io_out_0; // @[MUL.scala 124:19]
  wire  m_1997_io_out_1; // @[MUL.scala 124:19]
  wire  m_1998_io_x1; // @[MUL.scala 102:19]
  wire  m_1998_io_x2; // @[MUL.scala 102:19]
  wire  m_1998_io_x3; // @[MUL.scala 102:19]
  wire  m_1998_io_s; // @[MUL.scala 102:19]
  wire  m_1998_io_cout; // @[MUL.scala 102:19]
  wire  m_1999_io_in_0; // @[MUL.scala 124:19]
  wire  m_1999_io_in_1; // @[MUL.scala 124:19]
  wire  m_1999_io_out_0; // @[MUL.scala 124:19]
  wire  m_1999_io_out_1; // @[MUL.scala 124:19]
  wire  m_2000_io_x1; // @[MUL.scala 102:19]
  wire  m_2000_io_x2; // @[MUL.scala 102:19]
  wire  m_2000_io_x3; // @[MUL.scala 102:19]
  wire  m_2000_io_s; // @[MUL.scala 102:19]
  wire  m_2000_io_cout; // @[MUL.scala 102:19]
  wire  m_2001_io_in_0; // @[MUL.scala 124:19]
  wire  m_2001_io_in_1; // @[MUL.scala 124:19]
  wire  m_2001_io_out_0; // @[MUL.scala 124:19]
  wire  m_2001_io_out_1; // @[MUL.scala 124:19]
  wire  m_2002_io_x1; // @[MUL.scala 102:19]
  wire  m_2002_io_x2; // @[MUL.scala 102:19]
  wire  m_2002_io_x3; // @[MUL.scala 102:19]
  wire  m_2002_io_s; // @[MUL.scala 102:19]
  wire  m_2002_io_cout; // @[MUL.scala 102:19]
  wire  m_2003_io_x1; // @[MUL.scala 102:19]
  wire  m_2003_io_x2; // @[MUL.scala 102:19]
  wire  m_2003_io_x3; // @[MUL.scala 102:19]
  wire  m_2003_io_s; // @[MUL.scala 102:19]
  wire  m_2003_io_cout; // @[MUL.scala 102:19]
  wire  m_2004_io_x1; // @[MUL.scala 102:19]
  wire  m_2004_io_x2; // @[MUL.scala 102:19]
  wire  m_2004_io_x3; // @[MUL.scala 102:19]
  wire  m_2004_io_s; // @[MUL.scala 102:19]
  wire  m_2004_io_cout; // @[MUL.scala 102:19]
  wire  m_2005_io_x1; // @[MUL.scala 102:19]
  wire  m_2005_io_x2; // @[MUL.scala 102:19]
  wire  m_2005_io_x3; // @[MUL.scala 102:19]
  wire  m_2005_io_s; // @[MUL.scala 102:19]
  wire  m_2005_io_cout; // @[MUL.scala 102:19]
  wire  m_2006_io_x1; // @[MUL.scala 102:19]
  wire  m_2006_io_x2; // @[MUL.scala 102:19]
  wire  m_2006_io_x3; // @[MUL.scala 102:19]
  wire  m_2006_io_s; // @[MUL.scala 102:19]
  wire  m_2006_io_cout; // @[MUL.scala 102:19]
  wire  m_2007_io_x1; // @[MUL.scala 102:19]
  wire  m_2007_io_x2; // @[MUL.scala 102:19]
  wire  m_2007_io_x3; // @[MUL.scala 102:19]
  wire  m_2007_io_s; // @[MUL.scala 102:19]
  wire  m_2007_io_cout; // @[MUL.scala 102:19]
  wire  m_2008_io_x1; // @[MUL.scala 102:19]
  wire  m_2008_io_x2; // @[MUL.scala 102:19]
  wire  m_2008_io_x3; // @[MUL.scala 102:19]
  wire  m_2008_io_s; // @[MUL.scala 102:19]
  wire  m_2008_io_cout; // @[MUL.scala 102:19]
  wire  m_2009_io_x1; // @[MUL.scala 102:19]
  wire  m_2009_io_x2; // @[MUL.scala 102:19]
  wire  m_2009_io_x3; // @[MUL.scala 102:19]
  wire  m_2009_io_s; // @[MUL.scala 102:19]
  wire  m_2009_io_cout; // @[MUL.scala 102:19]
  wire  m_2010_io_x1; // @[MUL.scala 102:19]
  wire  m_2010_io_x2; // @[MUL.scala 102:19]
  wire  m_2010_io_x3; // @[MUL.scala 102:19]
  wire  m_2010_io_s; // @[MUL.scala 102:19]
  wire  m_2010_io_cout; // @[MUL.scala 102:19]
  wire  m_2011_io_x1; // @[MUL.scala 102:19]
  wire  m_2011_io_x2; // @[MUL.scala 102:19]
  wire  m_2011_io_x3; // @[MUL.scala 102:19]
  wire  m_2011_io_s; // @[MUL.scala 102:19]
  wire  m_2011_io_cout; // @[MUL.scala 102:19]
  wire  m_2012_io_x1; // @[MUL.scala 102:19]
  wire  m_2012_io_x2; // @[MUL.scala 102:19]
  wire  m_2012_io_x3; // @[MUL.scala 102:19]
  wire  m_2012_io_s; // @[MUL.scala 102:19]
  wire  m_2012_io_cout; // @[MUL.scala 102:19]
  wire  m_2013_io_x1; // @[MUL.scala 102:19]
  wire  m_2013_io_x2; // @[MUL.scala 102:19]
  wire  m_2013_io_x3; // @[MUL.scala 102:19]
  wire  m_2013_io_s; // @[MUL.scala 102:19]
  wire  m_2013_io_cout; // @[MUL.scala 102:19]
  wire  m_2014_io_x1; // @[MUL.scala 102:19]
  wire  m_2014_io_x2; // @[MUL.scala 102:19]
  wire  m_2014_io_x3; // @[MUL.scala 102:19]
  wire  m_2014_io_s; // @[MUL.scala 102:19]
  wire  m_2014_io_cout; // @[MUL.scala 102:19]
  wire  m_2015_io_x1; // @[MUL.scala 102:19]
  wire  m_2015_io_x2; // @[MUL.scala 102:19]
  wire  m_2015_io_x3; // @[MUL.scala 102:19]
  wire  m_2015_io_s; // @[MUL.scala 102:19]
  wire  m_2015_io_cout; // @[MUL.scala 102:19]
  wire  m_2016_io_x1; // @[MUL.scala 102:19]
  wire  m_2016_io_x2; // @[MUL.scala 102:19]
  wire  m_2016_io_x3; // @[MUL.scala 102:19]
  wire  m_2016_io_s; // @[MUL.scala 102:19]
  wire  m_2016_io_cout; // @[MUL.scala 102:19]
  wire  m_2017_io_x1; // @[MUL.scala 102:19]
  wire  m_2017_io_x2; // @[MUL.scala 102:19]
  wire  m_2017_io_x3; // @[MUL.scala 102:19]
  wire  m_2017_io_s; // @[MUL.scala 102:19]
  wire  m_2017_io_cout; // @[MUL.scala 102:19]
  wire  m_2018_io_x1; // @[MUL.scala 102:19]
  wire  m_2018_io_x2; // @[MUL.scala 102:19]
  wire  m_2018_io_x3; // @[MUL.scala 102:19]
  wire  m_2018_io_s; // @[MUL.scala 102:19]
  wire  m_2018_io_cout; // @[MUL.scala 102:19]
  wire  m_2019_io_x1; // @[MUL.scala 102:19]
  wire  m_2019_io_x2; // @[MUL.scala 102:19]
  wire  m_2019_io_x3; // @[MUL.scala 102:19]
  wire  m_2019_io_s; // @[MUL.scala 102:19]
  wire  m_2019_io_cout; // @[MUL.scala 102:19]
  wire  m_2020_io_x1; // @[MUL.scala 102:19]
  wire  m_2020_io_x2; // @[MUL.scala 102:19]
  wire  m_2020_io_x3; // @[MUL.scala 102:19]
  wire  m_2020_io_s; // @[MUL.scala 102:19]
  wire  m_2020_io_cout; // @[MUL.scala 102:19]
  wire  m_2021_io_x1; // @[MUL.scala 102:19]
  wire  m_2021_io_x2; // @[MUL.scala 102:19]
  wire  m_2021_io_x3; // @[MUL.scala 102:19]
  wire  m_2021_io_s; // @[MUL.scala 102:19]
  wire  m_2021_io_cout; // @[MUL.scala 102:19]
  wire  m_2022_io_x1; // @[MUL.scala 102:19]
  wire  m_2022_io_x2; // @[MUL.scala 102:19]
  wire  m_2022_io_x3; // @[MUL.scala 102:19]
  wire  m_2022_io_s; // @[MUL.scala 102:19]
  wire  m_2022_io_cout; // @[MUL.scala 102:19]
  wire  m_2023_io_x1; // @[MUL.scala 102:19]
  wire  m_2023_io_x2; // @[MUL.scala 102:19]
  wire  m_2023_io_x3; // @[MUL.scala 102:19]
  wire  m_2023_io_s; // @[MUL.scala 102:19]
  wire  m_2023_io_cout; // @[MUL.scala 102:19]
  wire  m_2024_io_x1; // @[MUL.scala 102:19]
  wire  m_2024_io_x2; // @[MUL.scala 102:19]
  wire  m_2024_io_x3; // @[MUL.scala 102:19]
  wire  m_2024_io_s; // @[MUL.scala 102:19]
  wire  m_2024_io_cout; // @[MUL.scala 102:19]
  wire  m_2025_io_x1; // @[MUL.scala 102:19]
  wire  m_2025_io_x2; // @[MUL.scala 102:19]
  wire  m_2025_io_x3; // @[MUL.scala 102:19]
  wire  m_2025_io_s; // @[MUL.scala 102:19]
  wire  m_2025_io_cout; // @[MUL.scala 102:19]
  wire  m_2026_io_x1; // @[MUL.scala 102:19]
  wire  m_2026_io_x2; // @[MUL.scala 102:19]
  wire  m_2026_io_x3; // @[MUL.scala 102:19]
  wire  m_2026_io_s; // @[MUL.scala 102:19]
  wire  m_2026_io_cout; // @[MUL.scala 102:19]
  wire  m_2027_io_x1; // @[MUL.scala 102:19]
  wire  m_2027_io_x2; // @[MUL.scala 102:19]
  wire  m_2027_io_x3; // @[MUL.scala 102:19]
  wire  m_2027_io_s; // @[MUL.scala 102:19]
  wire  m_2027_io_cout; // @[MUL.scala 102:19]
  wire  m_2028_io_x1; // @[MUL.scala 102:19]
  wire  m_2028_io_x2; // @[MUL.scala 102:19]
  wire  m_2028_io_x3; // @[MUL.scala 102:19]
  wire  m_2028_io_s; // @[MUL.scala 102:19]
  wire  m_2028_io_cout; // @[MUL.scala 102:19]
  wire  m_2029_io_x1; // @[MUL.scala 102:19]
  wire  m_2029_io_x2; // @[MUL.scala 102:19]
  wire  m_2029_io_x3; // @[MUL.scala 102:19]
  wire  m_2029_io_s; // @[MUL.scala 102:19]
  wire  m_2029_io_cout; // @[MUL.scala 102:19]
  wire  m_2030_io_x1; // @[MUL.scala 102:19]
  wire  m_2030_io_x2; // @[MUL.scala 102:19]
  wire  m_2030_io_x3; // @[MUL.scala 102:19]
  wire  m_2030_io_s; // @[MUL.scala 102:19]
  wire  m_2030_io_cout; // @[MUL.scala 102:19]
  wire  m_2031_io_x1; // @[MUL.scala 102:19]
  wire  m_2031_io_x2; // @[MUL.scala 102:19]
  wire  m_2031_io_x3; // @[MUL.scala 102:19]
  wire  m_2031_io_s; // @[MUL.scala 102:19]
  wire  m_2031_io_cout; // @[MUL.scala 102:19]
  wire  m_2032_io_x1; // @[MUL.scala 102:19]
  wire  m_2032_io_x2; // @[MUL.scala 102:19]
  wire  m_2032_io_x3; // @[MUL.scala 102:19]
  wire  m_2032_io_s; // @[MUL.scala 102:19]
  wire  m_2032_io_cout; // @[MUL.scala 102:19]
  wire  m_2033_io_x1; // @[MUL.scala 102:19]
  wire  m_2033_io_x2; // @[MUL.scala 102:19]
  wire  m_2033_io_x3; // @[MUL.scala 102:19]
  wire  m_2033_io_s; // @[MUL.scala 102:19]
  wire  m_2033_io_cout; // @[MUL.scala 102:19]
  wire  m_2034_io_x1; // @[MUL.scala 102:19]
  wire  m_2034_io_x2; // @[MUL.scala 102:19]
  wire  m_2034_io_x3; // @[MUL.scala 102:19]
  wire  m_2034_io_s; // @[MUL.scala 102:19]
  wire  m_2034_io_cout; // @[MUL.scala 102:19]
  wire  m_2035_io_x1; // @[MUL.scala 102:19]
  wire  m_2035_io_x2; // @[MUL.scala 102:19]
  wire  m_2035_io_x3; // @[MUL.scala 102:19]
  wire  m_2035_io_s; // @[MUL.scala 102:19]
  wire  m_2035_io_cout; // @[MUL.scala 102:19]
  wire  m_2036_io_x1; // @[MUL.scala 102:19]
  wire  m_2036_io_x2; // @[MUL.scala 102:19]
  wire  m_2036_io_x3; // @[MUL.scala 102:19]
  wire  m_2036_io_s; // @[MUL.scala 102:19]
  wire  m_2036_io_cout; // @[MUL.scala 102:19]
  wire  m_2037_io_x1; // @[MUL.scala 102:19]
  wire  m_2037_io_x2; // @[MUL.scala 102:19]
  wire  m_2037_io_x3; // @[MUL.scala 102:19]
  wire  m_2037_io_s; // @[MUL.scala 102:19]
  wire  m_2037_io_cout; // @[MUL.scala 102:19]
  wire  m_2038_io_x1; // @[MUL.scala 102:19]
  wire  m_2038_io_x2; // @[MUL.scala 102:19]
  wire  m_2038_io_x3; // @[MUL.scala 102:19]
  wire  m_2038_io_s; // @[MUL.scala 102:19]
  wire  m_2038_io_cout; // @[MUL.scala 102:19]
  wire  m_2039_io_x1; // @[MUL.scala 102:19]
  wire  m_2039_io_x2; // @[MUL.scala 102:19]
  wire  m_2039_io_x3; // @[MUL.scala 102:19]
  wire  m_2039_io_s; // @[MUL.scala 102:19]
  wire  m_2039_io_cout; // @[MUL.scala 102:19]
  wire  m_2040_io_x1; // @[MUL.scala 102:19]
  wire  m_2040_io_x2; // @[MUL.scala 102:19]
  wire  m_2040_io_x3; // @[MUL.scala 102:19]
  wire  m_2040_io_s; // @[MUL.scala 102:19]
  wire  m_2040_io_cout; // @[MUL.scala 102:19]
  wire  m_2041_io_x1; // @[MUL.scala 102:19]
  wire  m_2041_io_x2; // @[MUL.scala 102:19]
  wire  m_2041_io_x3; // @[MUL.scala 102:19]
  wire  m_2041_io_s; // @[MUL.scala 102:19]
  wire  m_2041_io_cout; // @[MUL.scala 102:19]
  wire  m_2042_io_x1; // @[MUL.scala 102:19]
  wire  m_2042_io_x2; // @[MUL.scala 102:19]
  wire  m_2042_io_x3; // @[MUL.scala 102:19]
  wire  m_2042_io_s; // @[MUL.scala 102:19]
  wire  m_2042_io_cout; // @[MUL.scala 102:19]
  wire  m_2043_io_x1; // @[MUL.scala 102:19]
  wire  m_2043_io_x2; // @[MUL.scala 102:19]
  wire  m_2043_io_x3; // @[MUL.scala 102:19]
  wire  m_2043_io_s; // @[MUL.scala 102:19]
  wire  m_2043_io_cout; // @[MUL.scala 102:19]
  wire  m_2044_io_x1; // @[MUL.scala 102:19]
  wire  m_2044_io_x2; // @[MUL.scala 102:19]
  wire  m_2044_io_x3; // @[MUL.scala 102:19]
  wire  m_2044_io_s; // @[MUL.scala 102:19]
  wire  m_2044_io_cout; // @[MUL.scala 102:19]
  wire  m_2045_io_x1; // @[MUL.scala 102:19]
  wire  m_2045_io_x2; // @[MUL.scala 102:19]
  wire  m_2045_io_x3; // @[MUL.scala 102:19]
  wire  m_2045_io_s; // @[MUL.scala 102:19]
  wire  m_2045_io_cout; // @[MUL.scala 102:19]
  wire  m_2046_io_x1; // @[MUL.scala 102:19]
  wire  m_2046_io_x2; // @[MUL.scala 102:19]
  wire  m_2046_io_x3; // @[MUL.scala 102:19]
  wire  m_2046_io_s; // @[MUL.scala 102:19]
  wire  m_2046_io_cout; // @[MUL.scala 102:19]
  wire  m_2047_io_x1; // @[MUL.scala 102:19]
  wire  m_2047_io_x2; // @[MUL.scala 102:19]
  wire  m_2047_io_x3; // @[MUL.scala 102:19]
  wire  m_2047_io_s; // @[MUL.scala 102:19]
  wire  m_2047_io_cout; // @[MUL.scala 102:19]
  wire  m_2048_io_x1; // @[MUL.scala 102:19]
  wire  m_2048_io_x2; // @[MUL.scala 102:19]
  wire  m_2048_io_x3; // @[MUL.scala 102:19]
  wire  m_2048_io_s; // @[MUL.scala 102:19]
  wire  m_2048_io_cout; // @[MUL.scala 102:19]
  wire  m_2049_io_x1; // @[MUL.scala 102:19]
  wire  m_2049_io_x2; // @[MUL.scala 102:19]
  wire  m_2049_io_x3; // @[MUL.scala 102:19]
  wire  m_2049_io_s; // @[MUL.scala 102:19]
  wire  m_2049_io_cout; // @[MUL.scala 102:19]
  wire  m_2050_io_x1; // @[MUL.scala 102:19]
  wire  m_2050_io_x2; // @[MUL.scala 102:19]
  wire  m_2050_io_x3; // @[MUL.scala 102:19]
  wire  m_2050_io_s; // @[MUL.scala 102:19]
  wire  m_2050_io_cout; // @[MUL.scala 102:19]
  wire  m_2051_io_x1; // @[MUL.scala 102:19]
  wire  m_2051_io_x2; // @[MUL.scala 102:19]
  wire  m_2051_io_x3; // @[MUL.scala 102:19]
  wire  m_2051_io_s; // @[MUL.scala 102:19]
  wire  m_2051_io_cout; // @[MUL.scala 102:19]
  wire  m_2052_io_x1; // @[MUL.scala 102:19]
  wire  m_2052_io_x2; // @[MUL.scala 102:19]
  wire  m_2052_io_x3; // @[MUL.scala 102:19]
  wire  m_2052_io_s; // @[MUL.scala 102:19]
  wire  m_2052_io_cout; // @[MUL.scala 102:19]
  wire  m_2053_io_x1; // @[MUL.scala 102:19]
  wire  m_2053_io_x2; // @[MUL.scala 102:19]
  wire  m_2053_io_x3; // @[MUL.scala 102:19]
  wire  m_2053_io_s; // @[MUL.scala 102:19]
  wire  m_2053_io_cout; // @[MUL.scala 102:19]
  wire  m_2054_io_x1; // @[MUL.scala 102:19]
  wire  m_2054_io_x2; // @[MUL.scala 102:19]
  wire  m_2054_io_x3; // @[MUL.scala 102:19]
  wire  m_2054_io_s; // @[MUL.scala 102:19]
  wire  m_2054_io_cout; // @[MUL.scala 102:19]
  wire  m_2055_io_x1; // @[MUL.scala 102:19]
  wire  m_2055_io_x2; // @[MUL.scala 102:19]
  wire  m_2055_io_x3; // @[MUL.scala 102:19]
  wire  m_2055_io_s; // @[MUL.scala 102:19]
  wire  m_2055_io_cout; // @[MUL.scala 102:19]
  wire  m_2056_io_x1; // @[MUL.scala 102:19]
  wire  m_2056_io_x2; // @[MUL.scala 102:19]
  wire  m_2056_io_x3; // @[MUL.scala 102:19]
  wire  m_2056_io_s; // @[MUL.scala 102:19]
  wire  m_2056_io_cout; // @[MUL.scala 102:19]
  wire  m_2057_io_x1; // @[MUL.scala 102:19]
  wire  m_2057_io_x2; // @[MUL.scala 102:19]
  wire  m_2057_io_x3; // @[MUL.scala 102:19]
  wire  m_2057_io_s; // @[MUL.scala 102:19]
  wire  m_2057_io_cout; // @[MUL.scala 102:19]
  wire  m_2058_io_x1; // @[MUL.scala 102:19]
  wire  m_2058_io_x2; // @[MUL.scala 102:19]
  wire  m_2058_io_x3; // @[MUL.scala 102:19]
  wire  m_2058_io_s; // @[MUL.scala 102:19]
  wire  m_2058_io_cout; // @[MUL.scala 102:19]
  wire  m_2059_io_x1; // @[MUL.scala 102:19]
  wire  m_2059_io_x2; // @[MUL.scala 102:19]
  wire  m_2059_io_x3; // @[MUL.scala 102:19]
  wire  m_2059_io_s; // @[MUL.scala 102:19]
  wire  m_2059_io_cout; // @[MUL.scala 102:19]
  wire  m_2060_io_x1; // @[MUL.scala 102:19]
  wire  m_2060_io_x2; // @[MUL.scala 102:19]
  wire  m_2060_io_x3; // @[MUL.scala 102:19]
  wire  m_2060_io_s; // @[MUL.scala 102:19]
  wire  m_2060_io_cout; // @[MUL.scala 102:19]
  wire  m_2061_io_x1; // @[MUL.scala 102:19]
  wire  m_2061_io_x2; // @[MUL.scala 102:19]
  wire  m_2061_io_x3; // @[MUL.scala 102:19]
  wire  m_2061_io_s; // @[MUL.scala 102:19]
  wire  m_2061_io_cout; // @[MUL.scala 102:19]
  wire  m_2062_io_x1; // @[MUL.scala 102:19]
  wire  m_2062_io_x2; // @[MUL.scala 102:19]
  wire  m_2062_io_x3; // @[MUL.scala 102:19]
  wire  m_2062_io_s; // @[MUL.scala 102:19]
  wire  m_2062_io_cout; // @[MUL.scala 102:19]
  wire  m_2063_io_x1; // @[MUL.scala 102:19]
  wire  m_2063_io_x2; // @[MUL.scala 102:19]
  wire  m_2063_io_x3; // @[MUL.scala 102:19]
  wire  m_2063_io_s; // @[MUL.scala 102:19]
  wire  m_2063_io_cout; // @[MUL.scala 102:19]
  wire  m_2064_io_x1; // @[MUL.scala 102:19]
  wire  m_2064_io_x2; // @[MUL.scala 102:19]
  wire  m_2064_io_x3; // @[MUL.scala 102:19]
  wire  m_2064_io_s; // @[MUL.scala 102:19]
  wire  m_2064_io_cout; // @[MUL.scala 102:19]
  wire  m_2065_io_x1; // @[MUL.scala 102:19]
  wire  m_2065_io_x2; // @[MUL.scala 102:19]
  wire  m_2065_io_x3; // @[MUL.scala 102:19]
  wire  m_2065_io_s; // @[MUL.scala 102:19]
  wire  m_2065_io_cout; // @[MUL.scala 102:19]
  wire  m_2066_io_x1; // @[MUL.scala 102:19]
  wire  m_2066_io_x2; // @[MUL.scala 102:19]
  wire  m_2066_io_x3; // @[MUL.scala 102:19]
  wire  m_2066_io_s; // @[MUL.scala 102:19]
  wire  m_2066_io_cout; // @[MUL.scala 102:19]
  wire  m_2067_io_x1; // @[MUL.scala 102:19]
  wire  m_2067_io_x2; // @[MUL.scala 102:19]
  wire  m_2067_io_x3; // @[MUL.scala 102:19]
  wire  m_2067_io_s; // @[MUL.scala 102:19]
  wire  m_2067_io_cout; // @[MUL.scala 102:19]
  wire  m_2068_io_x1; // @[MUL.scala 102:19]
  wire  m_2068_io_x2; // @[MUL.scala 102:19]
  wire  m_2068_io_x3; // @[MUL.scala 102:19]
  wire  m_2068_io_s; // @[MUL.scala 102:19]
  wire  m_2068_io_cout; // @[MUL.scala 102:19]
  wire  m_2069_io_x1; // @[MUL.scala 102:19]
  wire  m_2069_io_x2; // @[MUL.scala 102:19]
  wire  m_2069_io_x3; // @[MUL.scala 102:19]
  wire  m_2069_io_s; // @[MUL.scala 102:19]
  wire  m_2069_io_cout; // @[MUL.scala 102:19]
  wire  m_2070_io_x1; // @[MUL.scala 102:19]
  wire  m_2070_io_x2; // @[MUL.scala 102:19]
  wire  m_2070_io_x3; // @[MUL.scala 102:19]
  wire  m_2070_io_s; // @[MUL.scala 102:19]
  wire  m_2070_io_cout; // @[MUL.scala 102:19]
  wire  m_2071_io_x1; // @[MUL.scala 102:19]
  wire  m_2071_io_x2; // @[MUL.scala 102:19]
  wire  m_2071_io_x3; // @[MUL.scala 102:19]
  wire  m_2071_io_s; // @[MUL.scala 102:19]
  wire  m_2071_io_cout; // @[MUL.scala 102:19]
  wire  m_2072_io_x1; // @[MUL.scala 102:19]
  wire  m_2072_io_x2; // @[MUL.scala 102:19]
  wire  m_2072_io_x3; // @[MUL.scala 102:19]
  wire  m_2072_io_s; // @[MUL.scala 102:19]
  wire  m_2072_io_cout; // @[MUL.scala 102:19]
  wire  m_2073_io_x1; // @[MUL.scala 102:19]
  wire  m_2073_io_x2; // @[MUL.scala 102:19]
  wire  m_2073_io_x3; // @[MUL.scala 102:19]
  wire  m_2073_io_s; // @[MUL.scala 102:19]
  wire  m_2073_io_cout; // @[MUL.scala 102:19]
  wire  m_2074_io_x1; // @[MUL.scala 102:19]
  wire  m_2074_io_x2; // @[MUL.scala 102:19]
  wire  m_2074_io_x3; // @[MUL.scala 102:19]
  wire  m_2074_io_s; // @[MUL.scala 102:19]
  wire  m_2074_io_cout; // @[MUL.scala 102:19]
  wire  m_2075_io_x1; // @[MUL.scala 102:19]
  wire  m_2075_io_x2; // @[MUL.scala 102:19]
  wire  m_2075_io_x3; // @[MUL.scala 102:19]
  wire  m_2075_io_s; // @[MUL.scala 102:19]
  wire  m_2075_io_cout; // @[MUL.scala 102:19]
  wire  m_2076_io_x1; // @[MUL.scala 102:19]
  wire  m_2076_io_x2; // @[MUL.scala 102:19]
  wire  m_2076_io_x3; // @[MUL.scala 102:19]
  wire  m_2076_io_s; // @[MUL.scala 102:19]
  wire  m_2076_io_cout; // @[MUL.scala 102:19]
  wire  m_2077_io_x1; // @[MUL.scala 102:19]
  wire  m_2077_io_x2; // @[MUL.scala 102:19]
  wire  m_2077_io_x3; // @[MUL.scala 102:19]
  wire  m_2077_io_s; // @[MUL.scala 102:19]
  wire  m_2077_io_cout; // @[MUL.scala 102:19]
  wire  m_2078_io_x1; // @[MUL.scala 102:19]
  wire  m_2078_io_x2; // @[MUL.scala 102:19]
  wire  m_2078_io_x3; // @[MUL.scala 102:19]
  wire  m_2078_io_s; // @[MUL.scala 102:19]
  wire  m_2078_io_cout; // @[MUL.scala 102:19]
  wire  m_2079_io_x1; // @[MUL.scala 102:19]
  wire  m_2079_io_x2; // @[MUL.scala 102:19]
  wire  m_2079_io_x3; // @[MUL.scala 102:19]
  wire  m_2079_io_s; // @[MUL.scala 102:19]
  wire  m_2079_io_cout; // @[MUL.scala 102:19]
  wire  m_2080_io_x1; // @[MUL.scala 102:19]
  wire  m_2080_io_x2; // @[MUL.scala 102:19]
  wire  m_2080_io_x3; // @[MUL.scala 102:19]
  wire  m_2080_io_s; // @[MUL.scala 102:19]
  wire  m_2080_io_cout; // @[MUL.scala 102:19]
  wire  m_2081_io_x1; // @[MUL.scala 102:19]
  wire  m_2081_io_x2; // @[MUL.scala 102:19]
  wire  m_2081_io_x3; // @[MUL.scala 102:19]
  wire  m_2081_io_s; // @[MUL.scala 102:19]
  wire  m_2081_io_cout; // @[MUL.scala 102:19]
  wire  m_2082_io_x1; // @[MUL.scala 102:19]
  wire  m_2082_io_x2; // @[MUL.scala 102:19]
  wire  m_2082_io_x3; // @[MUL.scala 102:19]
  wire  m_2082_io_s; // @[MUL.scala 102:19]
  wire  m_2082_io_cout; // @[MUL.scala 102:19]
  wire  m_2083_io_x1; // @[MUL.scala 102:19]
  wire  m_2083_io_x2; // @[MUL.scala 102:19]
  wire  m_2083_io_x3; // @[MUL.scala 102:19]
  wire  m_2083_io_s; // @[MUL.scala 102:19]
  wire  m_2083_io_cout; // @[MUL.scala 102:19]
  wire  m_2084_io_x1; // @[MUL.scala 102:19]
  wire  m_2084_io_x2; // @[MUL.scala 102:19]
  wire  m_2084_io_x3; // @[MUL.scala 102:19]
  wire  m_2084_io_s; // @[MUL.scala 102:19]
  wire  m_2084_io_cout; // @[MUL.scala 102:19]
  wire  m_2085_io_x1; // @[MUL.scala 102:19]
  wire  m_2085_io_x2; // @[MUL.scala 102:19]
  wire  m_2085_io_x3; // @[MUL.scala 102:19]
  wire  m_2085_io_s; // @[MUL.scala 102:19]
  wire  m_2085_io_cout; // @[MUL.scala 102:19]
  wire  m_2086_io_x1; // @[MUL.scala 102:19]
  wire  m_2086_io_x2; // @[MUL.scala 102:19]
  wire  m_2086_io_x3; // @[MUL.scala 102:19]
  wire  m_2086_io_s; // @[MUL.scala 102:19]
  wire  m_2086_io_cout; // @[MUL.scala 102:19]
  wire  m_2087_io_x1; // @[MUL.scala 102:19]
  wire  m_2087_io_x2; // @[MUL.scala 102:19]
  wire  m_2087_io_x3; // @[MUL.scala 102:19]
  wire  m_2087_io_s; // @[MUL.scala 102:19]
  wire  m_2087_io_cout; // @[MUL.scala 102:19]
  wire  m_2088_io_x1; // @[MUL.scala 102:19]
  wire  m_2088_io_x2; // @[MUL.scala 102:19]
  wire  m_2088_io_x3; // @[MUL.scala 102:19]
  wire  m_2088_io_s; // @[MUL.scala 102:19]
  wire  m_2088_io_cout; // @[MUL.scala 102:19]
  wire  m_2089_io_x1; // @[MUL.scala 102:19]
  wire  m_2089_io_x2; // @[MUL.scala 102:19]
  wire  m_2089_io_x3; // @[MUL.scala 102:19]
  wire  m_2089_io_s; // @[MUL.scala 102:19]
  wire  m_2089_io_cout; // @[MUL.scala 102:19]
  wire  m_2090_io_x1; // @[MUL.scala 102:19]
  wire  m_2090_io_x2; // @[MUL.scala 102:19]
  wire  m_2090_io_x3; // @[MUL.scala 102:19]
  wire  m_2090_io_s; // @[MUL.scala 102:19]
  wire  m_2090_io_cout; // @[MUL.scala 102:19]
  wire  m_2091_io_x1; // @[MUL.scala 102:19]
  wire  m_2091_io_x2; // @[MUL.scala 102:19]
  wire  m_2091_io_x3; // @[MUL.scala 102:19]
  wire  m_2091_io_s; // @[MUL.scala 102:19]
  wire  m_2091_io_cout; // @[MUL.scala 102:19]
  wire  m_2092_io_x1; // @[MUL.scala 102:19]
  wire  m_2092_io_x2; // @[MUL.scala 102:19]
  wire  m_2092_io_x3; // @[MUL.scala 102:19]
  wire  m_2092_io_s; // @[MUL.scala 102:19]
  wire  m_2092_io_cout; // @[MUL.scala 102:19]
  wire  m_2093_io_x1; // @[MUL.scala 102:19]
  wire  m_2093_io_x2; // @[MUL.scala 102:19]
  wire  m_2093_io_x3; // @[MUL.scala 102:19]
  wire  m_2093_io_s; // @[MUL.scala 102:19]
  wire  m_2093_io_cout; // @[MUL.scala 102:19]
  wire  m_2094_io_x1; // @[MUL.scala 102:19]
  wire  m_2094_io_x2; // @[MUL.scala 102:19]
  wire  m_2094_io_x3; // @[MUL.scala 102:19]
  wire  m_2094_io_s; // @[MUL.scala 102:19]
  wire  m_2094_io_cout; // @[MUL.scala 102:19]
  wire  m_2095_io_in_0; // @[MUL.scala 124:19]
  wire  m_2095_io_in_1; // @[MUL.scala 124:19]
  wire  m_2095_io_out_0; // @[MUL.scala 124:19]
  wire  m_2095_io_out_1; // @[MUL.scala 124:19]
  wire  m_2096_io_x1; // @[MUL.scala 102:19]
  wire  m_2096_io_x2; // @[MUL.scala 102:19]
  wire  m_2096_io_x3; // @[MUL.scala 102:19]
  wire  m_2096_io_s; // @[MUL.scala 102:19]
  wire  m_2096_io_cout; // @[MUL.scala 102:19]
  wire  m_2097_io_in_0; // @[MUL.scala 124:19]
  wire  m_2097_io_in_1; // @[MUL.scala 124:19]
  wire  m_2097_io_out_0; // @[MUL.scala 124:19]
  wire  m_2097_io_out_1; // @[MUL.scala 124:19]
  wire  m_2098_io_x1; // @[MUL.scala 102:19]
  wire  m_2098_io_x2; // @[MUL.scala 102:19]
  wire  m_2098_io_x3; // @[MUL.scala 102:19]
  wire  m_2098_io_s; // @[MUL.scala 102:19]
  wire  m_2098_io_cout; // @[MUL.scala 102:19]
  wire  m_2099_io_in_0; // @[MUL.scala 124:19]
  wire  m_2099_io_in_1; // @[MUL.scala 124:19]
  wire  m_2099_io_out_0; // @[MUL.scala 124:19]
  wire  m_2099_io_out_1; // @[MUL.scala 124:19]
  wire  m_2100_io_x1; // @[MUL.scala 102:19]
  wire  m_2100_io_x2; // @[MUL.scala 102:19]
  wire  m_2100_io_x3; // @[MUL.scala 102:19]
  wire  m_2100_io_s; // @[MUL.scala 102:19]
  wire  m_2100_io_cout; // @[MUL.scala 102:19]
  wire  m_2101_io_in_0; // @[MUL.scala 124:19]
  wire  m_2101_io_in_1; // @[MUL.scala 124:19]
  wire  m_2101_io_out_0; // @[MUL.scala 124:19]
  wire  m_2101_io_out_1; // @[MUL.scala 124:19]
  wire  m_2102_io_x1; // @[MUL.scala 102:19]
  wire  m_2102_io_x2; // @[MUL.scala 102:19]
  wire  m_2102_io_x3; // @[MUL.scala 102:19]
  wire  m_2102_io_s; // @[MUL.scala 102:19]
  wire  m_2102_io_cout; // @[MUL.scala 102:19]
  wire  m_2103_io_in_0; // @[MUL.scala 124:19]
  wire  m_2103_io_in_1; // @[MUL.scala 124:19]
  wire  m_2103_io_out_0; // @[MUL.scala 124:19]
  wire  m_2103_io_out_1; // @[MUL.scala 124:19]
  wire  m_2104_io_x1; // @[MUL.scala 102:19]
  wire  m_2104_io_x2; // @[MUL.scala 102:19]
  wire  m_2104_io_x3; // @[MUL.scala 102:19]
  wire  m_2104_io_s; // @[MUL.scala 102:19]
  wire  m_2104_io_cout; // @[MUL.scala 102:19]
  wire  m_2105_io_x1; // @[MUL.scala 102:19]
  wire  m_2105_io_x2; // @[MUL.scala 102:19]
  wire  m_2105_io_x3; // @[MUL.scala 102:19]
  wire  m_2105_io_s; // @[MUL.scala 102:19]
  wire  m_2105_io_cout; // @[MUL.scala 102:19]
  wire  m_2106_io_x1; // @[MUL.scala 102:19]
  wire  m_2106_io_x2; // @[MUL.scala 102:19]
  wire  m_2106_io_x3; // @[MUL.scala 102:19]
  wire  m_2106_io_s; // @[MUL.scala 102:19]
  wire  m_2106_io_cout; // @[MUL.scala 102:19]
  wire  m_2107_io_x1; // @[MUL.scala 102:19]
  wire  m_2107_io_x2; // @[MUL.scala 102:19]
  wire  m_2107_io_x3; // @[MUL.scala 102:19]
  wire  m_2107_io_s; // @[MUL.scala 102:19]
  wire  m_2107_io_cout; // @[MUL.scala 102:19]
  wire  m_2108_io_x1; // @[MUL.scala 102:19]
  wire  m_2108_io_x2; // @[MUL.scala 102:19]
  wire  m_2108_io_x3; // @[MUL.scala 102:19]
  wire  m_2108_io_s; // @[MUL.scala 102:19]
  wire  m_2108_io_cout; // @[MUL.scala 102:19]
  wire  m_2109_io_x1; // @[MUL.scala 102:19]
  wire  m_2109_io_x2; // @[MUL.scala 102:19]
  wire  m_2109_io_x3; // @[MUL.scala 102:19]
  wire  m_2109_io_s; // @[MUL.scala 102:19]
  wire  m_2109_io_cout; // @[MUL.scala 102:19]
  wire  m_2110_io_x1; // @[MUL.scala 102:19]
  wire  m_2110_io_x2; // @[MUL.scala 102:19]
  wire  m_2110_io_x3; // @[MUL.scala 102:19]
  wire  m_2110_io_s; // @[MUL.scala 102:19]
  wire  m_2110_io_cout; // @[MUL.scala 102:19]
  wire  m_2111_io_x1; // @[MUL.scala 102:19]
  wire  m_2111_io_x2; // @[MUL.scala 102:19]
  wire  m_2111_io_x3; // @[MUL.scala 102:19]
  wire  m_2111_io_s; // @[MUL.scala 102:19]
  wire  m_2111_io_cout; // @[MUL.scala 102:19]
  wire  m_2112_io_x1; // @[MUL.scala 102:19]
  wire  m_2112_io_x2; // @[MUL.scala 102:19]
  wire  m_2112_io_x3; // @[MUL.scala 102:19]
  wire  m_2112_io_s; // @[MUL.scala 102:19]
  wire  m_2112_io_cout; // @[MUL.scala 102:19]
  wire  m_2113_io_x1; // @[MUL.scala 102:19]
  wire  m_2113_io_x2; // @[MUL.scala 102:19]
  wire  m_2113_io_x3; // @[MUL.scala 102:19]
  wire  m_2113_io_s; // @[MUL.scala 102:19]
  wire  m_2113_io_cout; // @[MUL.scala 102:19]
  wire  m_2114_io_x1; // @[MUL.scala 102:19]
  wire  m_2114_io_x2; // @[MUL.scala 102:19]
  wire  m_2114_io_x3; // @[MUL.scala 102:19]
  wire  m_2114_io_s; // @[MUL.scala 102:19]
  wire  m_2114_io_cout; // @[MUL.scala 102:19]
  wire  m_2115_io_x1; // @[MUL.scala 102:19]
  wire  m_2115_io_x2; // @[MUL.scala 102:19]
  wire  m_2115_io_x3; // @[MUL.scala 102:19]
  wire  m_2115_io_s; // @[MUL.scala 102:19]
  wire  m_2115_io_cout; // @[MUL.scala 102:19]
  wire  m_2116_io_x1; // @[MUL.scala 102:19]
  wire  m_2116_io_x2; // @[MUL.scala 102:19]
  wire  m_2116_io_x3; // @[MUL.scala 102:19]
  wire  m_2116_io_s; // @[MUL.scala 102:19]
  wire  m_2116_io_cout; // @[MUL.scala 102:19]
  wire  m_2117_io_x1; // @[MUL.scala 102:19]
  wire  m_2117_io_x2; // @[MUL.scala 102:19]
  wire  m_2117_io_x3; // @[MUL.scala 102:19]
  wire  m_2117_io_s; // @[MUL.scala 102:19]
  wire  m_2117_io_cout; // @[MUL.scala 102:19]
  wire  m_2118_io_x1; // @[MUL.scala 102:19]
  wire  m_2118_io_x2; // @[MUL.scala 102:19]
  wire  m_2118_io_x3; // @[MUL.scala 102:19]
  wire  m_2118_io_s; // @[MUL.scala 102:19]
  wire  m_2118_io_cout; // @[MUL.scala 102:19]
  wire  m_2119_io_x1; // @[MUL.scala 102:19]
  wire  m_2119_io_x2; // @[MUL.scala 102:19]
  wire  m_2119_io_x3; // @[MUL.scala 102:19]
  wire  m_2119_io_s; // @[MUL.scala 102:19]
  wire  m_2119_io_cout; // @[MUL.scala 102:19]
  wire  m_2120_io_x1; // @[MUL.scala 102:19]
  wire  m_2120_io_x2; // @[MUL.scala 102:19]
  wire  m_2120_io_x3; // @[MUL.scala 102:19]
  wire  m_2120_io_s; // @[MUL.scala 102:19]
  wire  m_2120_io_cout; // @[MUL.scala 102:19]
  wire  m_2121_io_x1; // @[MUL.scala 102:19]
  wire  m_2121_io_x2; // @[MUL.scala 102:19]
  wire  m_2121_io_x3; // @[MUL.scala 102:19]
  wire  m_2121_io_s; // @[MUL.scala 102:19]
  wire  m_2121_io_cout; // @[MUL.scala 102:19]
  wire  m_2122_io_x1; // @[MUL.scala 102:19]
  wire  m_2122_io_x2; // @[MUL.scala 102:19]
  wire  m_2122_io_x3; // @[MUL.scala 102:19]
  wire  m_2122_io_s; // @[MUL.scala 102:19]
  wire  m_2122_io_cout; // @[MUL.scala 102:19]
  wire  m_2123_io_in_0; // @[MUL.scala 124:19]
  wire  m_2123_io_in_1; // @[MUL.scala 124:19]
  wire  m_2123_io_out_0; // @[MUL.scala 124:19]
  wire  m_2123_io_out_1; // @[MUL.scala 124:19]
  wire  m_2124_io_in_0; // @[MUL.scala 124:19]
  wire  m_2124_io_in_1; // @[MUL.scala 124:19]
  wire  m_2124_io_out_0; // @[MUL.scala 124:19]
  wire  m_2124_io_out_1; // @[MUL.scala 124:19]
  wire  m_2125_io_in_0; // @[MUL.scala 124:19]
  wire  m_2125_io_in_1; // @[MUL.scala 124:19]
  wire  m_2125_io_out_0; // @[MUL.scala 124:19]
  wire  m_2125_io_out_1; // @[MUL.scala 124:19]
  wire  m_2126_io_in_0; // @[MUL.scala 124:19]
  wire  m_2126_io_in_1; // @[MUL.scala 124:19]
  wire  m_2126_io_out_0; // @[MUL.scala 124:19]
  wire  m_2126_io_out_1; // @[MUL.scala 124:19]
  wire  m_2127_io_in_0; // @[MUL.scala 124:19]
  wire  m_2127_io_in_1; // @[MUL.scala 124:19]
  wire  m_2127_io_out_0; // @[MUL.scala 124:19]
  wire  m_2127_io_out_1; // @[MUL.scala 124:19]
  wire  m_2128_io_in_0; // @[MUL.scala 124:19]
  wire  m_2128_io_in_1; // @[MUL.scala 124:19]
  wire  m_2128_io_out_0; // @[MUL.scala 124:19]
  wire  m_2128_io_out_1; // @[MUL.scala 124:19]
  wire  m_2129_io_in_0; // @[MUL.scala 124:19]
  wire  m_2129_io_in_1; // @[MUL.scala 124:19]
  wire  m_2129_io_out_0; // @[MUL.scala 124:19]
  wire  m_2129_io_out_1; // @[MUL.scala 124:19]
  wire  m_2130_io_in_0; // @[MUL.scala 124:19]
  wire  m_2130_io_in_1; // @[MUL.scala 124:19]
  wire  m_2130_io_out_0; // @[MUL.scala 124:19]
  wire  m_2130_io_out_1; // @[MUL.scala 124:19]
  wire  m_2131_io_in_0; // @[MUL.scala 124:19]
  wire  m_2131_io_in_1; // @[MUL.scala 124:19]
  wire  m_2131_io_out_0; // @[MUL.scala 124:19]
  wire  m_2131_io_out_1; // @[MUL.scala 124:19]
  wire  m_2132_io_in_0; // @[MUL.scala 124:19]
  wire  m_2132_io_in_1; // @[MUL.scala 124:19]
  wire  m_2132_io_out_0; // @[MUL.scala 124:19]
  wire  m_2132_io_out_1; // @[MUL.scala 124:19]
  wire  m_2133_io_in_0; // @[MUL.scala 124:19]
  wire  m_2133_io_in_1; // @[MUL.scala 124:19]
  wire  m_2133_io_out_0; // @[MUL.scala 124:19]
  wire  m_2133_io_out_1; // @[MUL.scala 124:19]
  wire  m_2134_io_in_0; // @[MUL.scala 124:19]
  wire  m_2134_io_in_1; // @[MUL.scala 124:19]
  wire  m_2134_io_out_0; // @[MUL.scala 124:19]
  wire  m_2134_io_out_1; // @[MUL.scala 124:19]
  wire  m_2135_io_in_0; // @[MUL.scala 124:19]
  wire  m_2135_io_in_1; // @[MUL.scala 124:19]
  wire  m_2135_io_out_0; // @[MUL.scala 124:19]
  wire  m_2135_io_out_1; // @[MUL.scala 124:19]
  wire  m_2136_io_in_0; // @[MUL.scala 124:19]
  wire  m_2136_io_in_1; // @[MUL.scala 124:19]
  wire  m_2136_io_out_0; // @[MUL.scala 124:19]
  wire  m_2136_io_out_1; // @[MUL.scala 124:19]
  wire  m_2137_io_in_0; // @[MUL.scala 124:19]
  wire  m_2137_io_in_1; // @[MUL.scala 124:19]
  wire  m_2137_io_out_0; // @[MUL.scala 124:19]
  wire  m_2137_io_out_1; // @[MUL.scala 124:19]
  wire  m_2138_io_in_0; // @[MUL.scala 124:19]
  wire  m_2138_io_in_1; // @[MUL.scala 124:19]
  wire  m_2138_io_out_0; // @[MUL.scala 124:19]
  wire  m_2138_io_out_1; // @[MUL.scala 124:19]
  wire  m_2139_io_in_0; // @[MUL.scala 124:19]
  wire  m_2139_io_in_1; // @[MUL.scala 124:19]
  wire  m_2139_io_out_0; // @[MUL.scala 124:19]
  wire  m_2139_io_out_1; // @[MUL.scala 124:19]
  wire  m_2140_io_in_0; // @[MUL.scala 124:19]
  wire  m_2140_io_in_1; // @[MUL.scala 124:19]
  wire  m_2140_io_out_0; // @[MUL.scala 124:19]
  wire  m_2140_io_out_1; // @[MUL.scala 124:19]
  wire  m_2141_io_in_0; // @[MUL.scala 124:19]
  wire  m_2141_io_in_1; // @[MUL.scala 124:19]
  wire  m_2141_io_out_0; // @[MUL.scala 124:19]
  wire  m_2141_io_out_1; // @[MUL.scala 124:19]
  wire  m_2142_io_in_0; // @[MUL.scala 124:19]
  wire  m_2142_io_in_1; // @[MUL.scala 124:19]
  wire  m_2142_io_out_0; // @[MUL.scala 124:19]
  wire  m_2142_io_out_1; // @[MUL.scala 124:19]
  wire  m_2143_io_in_0; // @[MUL.scala 124:19]
  wire  m_2143_io_in_1; // @[MUL.scala 124:19]
  wire  m_2143_io_out_0; // @[MUL.scala 124:19]
  wire  m_2143_io_out_1; // @[MUL.scala 124:19]
  wire  m_2144_io_in_0; // @[MUL.scala 124:19]
  wire  m_2144_io_in_1; // @[MUL.scala 124:19]
  wire  m_2144_io_out_0; // @[MUL.scala 124:19]
  wire  m_2144_io_out_1; // @[MUL.scala 124:19]
  wire  m_2145_io_in_0; // @[MUL.scala 124:19]
  wire  m_2145_io_in_1; // @[MUL.scala 124:19]
  wire  m_2145_io_out_0; // @[MUL.scala 124:19]
  wire  m_2145_io_out_1; // @[MUL.scala 124:19]
  wire  m_2146_io_in_0; // @[MUL.scala 124:19]
  wire  m_2146_io_in_1; // @[MUL.scala 124:19]
  wire  m_2146_io_out_0; // @[MUL.scala 124:19]
  wire  m_2146_io_out_1; // @[MUL.scala 124:19]
  wire  m_2147_io_in_0; // @[MUL.scala 124:19]
  wire  m_2147_io_in_1; // @[MUL.scala 124:19]
  wire  m_2147_io_out_0; // @[MUL.scala 124:19]
  wire  m_2147_io_out_1; // @[MUL.scala 124:19]
  wire  m_2148_io_in_0; // @[MUL.scala 124:19]
  wire  m_2148_io_in_1; // @[MUL.scala 124:19]
  wire  m_2148_io_out_0; // @[MUL.scala 124:19]
  wire  m_2148_io_out_1; // @[MUL.scala 124:19]
  wire  m_2149_io_in_0; // @[MUL.scala 124:19]
  wire  m_2149_io_in_1; // @[MUL.scala 124:19]
  wire  m_2149_io_out_0; // @[MUL.scala 124:19]
  wire  m_2149_io_out_1; // @[MUL.scala 124:19]
  wire  m_2150_io_in_0; // @[MUL.scala 124:19]
  wire  m_2150_io_in_1; // @[MUL.scala 124:19]
  wire  m_2150_io_out_0; // @[MUL.scala 124:19]
  wire  m_2150_io_out_1; // @[MUL.scala 124:19]
  wire  m_2151_io_in_0; // @[MUL.scala 124:19]
  wire  m_2151_io_in_1; // @[MUL.scala 124:19]
  wire  m_2151_io_out_0; // @[MUL.scala 124:19]
  wire  m_2151_io_out_1; // @[MUL.scala 124:19]
  wire  m_2152_io_in_0; // @[MUL.scala 124:19]
  wire  m_2152_io_in_1; // @[MUL.scala 124:19]
  wire  m_2152_io_out_0; // @[MUL.scala 124:19]
  wire  m_2152_io_out_1; // @[MUL.scala 124:19]
  wire  m_2153_io_in_0; // @[MUL.scala 124:19]
  wire  m_2153_io_in_1; // @[MUL.scala 124:19]
  wire  m_2153_io_out_0; // @[MUL.scala 124:19]
  wire  m_2153_io_out_1; // @[MUL.scala 124:19]
  wire  m_2154_io_in_0; // @[MUL.scala 124:19]
  wire  m_2154_io_in_1; // @[MUL.scala 124:19]
  wire  m_2154_io_out_0; // @[MUL.scala 124:19]
  wire  m_2154_io_out_1; // @[MUL.scala 124:19]
  wire  m_2155_io_in_0; // @[MUL.scala 124:19]
  wire  m_2155_io_in_1; // @[MUL.scala 124:19]
  wire  m_2155_io_out_0; // @[MUL.scala 124:19]
  wire  m_2155_io_out_1; // @[MUL.scala 124:19]
  wire  m_2156_io_in_0; // @[MUL.scala 124:19]
  wire  m_2156_io_in_1; // @[MUL.scala 124:19]
  wire  m_2156_io_out_0; // @[MUL.scala 124:19]
  wire  m_2156_io_out_1; // @[MUL.scala 124:19]
  wire  m_2157_io_in_0; // @[MUL.scala 124:19]
  wire  m_2157_io_in_1; // @[MUL.scala 124:19]
  wire  m_2157_io_out_0; // @[MUL.scala 124:19]
  wire  m_2157_io_out_1; // @[MUL.scala 124:19]
  wire  m_2158_io_in_0; // @[MUL.scala 124:19]
  wire  m_2158_io_in_1; // @[MUL.scala 124:19]
  wire  m_2158_io_out_0; // @[MUL.scala 124:19]
  wire  m_2158_io_out_1; // @[MUL.scala 124:19]
  wire  m_2159_io_in_0; // @[MUL.scala 124:19]
  wire  m_2159_io_in_1; // @[MUL.scala 124:19]
  wire  m_2159_io_out_0; // @[MUL.scala 124:19]
  wire  m_2159_io_out_1; // @[MUL.scala 124:19]
  wire  m_2160_io_x1; // @[MUL.scala 102:19]
  wire  m_2160_io_x2; // @[MUL.scala 102:19]
  wire  m_2160_io_x3; // @[MUL.scala 102:19]
  wire  m_2160_io_s; // @[MUL.scala 102:19]
  wire  m_2160_io_cout; // @[MUL.scala 102:19]
  wire  m_2161_io_x1; // @[MUL.scala 102:19]
  wire  m_2161_io_x2; // @[MUL.scala 102:19]
  wire  m_2161_io_x3; // @[MUL.scala 102:19]
  wire  m_2161_io_s; // @[MUL.scala 102:19]
  wire  m_2161_io_cout; // @[MUL.scala 102:19]
  wire  m_2162_io_x1; // @[MUL.scala 102:19]
  wire  m_2162_io_x2; // @[MUL.scala 102:19]
  wire  m_2162_io_x3; // @[MUL.scala 102:19]
  wire  m_2162_io_s; // @[MUL.scala 102:19]
  wire  m_2162_io_cout; // @[MUL.scala 102:19]
  wire  m_2163_io_x1; // @[MUL.scala 102:19]
  wire  m_2163_io_x2; // @[MUL.scala 102:19]
  wire  m_2163_io_x3; // @[MUL.scala 102:19]
  wire  m_2163_io_s; // @[MUL.scala 102:19]
  wire  m_2163_io_cout; // @[MUL.scala 102:19]
  wire  m_2164_io_x1; // @[MUL.scala 102:19]
  wire  m_2164_io_x2; // @[MUL.scala 102:19]
  wire  m_2164_io_x3; // @[MUL.scala 102:19]
  wire  m_2164_io_s; // @[MUL.scala 102:19]
  wire  m_2164_io_cout; // @[MUL.scala 102:19]
  wire  m_2165_io_x1; // @[MUL.scala 102:19]
  wire  m_2165_io_x2; // @[MUL.scala 102:19]
  wire  m_2165_io_x3; // @[MUL.scala 102:19]
  wire  m_2165_io_s; // @[MUL.scala 102:19]
  wire  m_2165_io_cout; // @[MUL.scala 102:19]
  wire  m_2166_io_x1; // @[MUL.scala 102:19]
  wire  m_2166_io_x2; // @[MUL.scala 102:19]
  wire  m_2166_io_x3; // @[MUL.scala 102:19]
  wire  m_2166_io_s; // @[MUL.scala 102:19]
  wire  m_2166_io_cout; // @[MUL.scala 102:19]
  wire  m_2167_io_x1; // @[MUL.scala 102:19]
  wire  m_2167_io_x2; // @[MUL.scala 102:19]
  wire  m_2167_io_x3; // @[MUL.scala 102:19]
  wire  m_2167_io_s; // @[MUL.scala 102:19]
  wire  m_2167_io_cout; // @[MUL.scala 102:19]
  wire  m_2168_io_x1; // @[MUL.scala 102:19]
  wire  m_2168_io_x2; // @[MUL.scala 102:19]
  wire  m_2168_io_x3; // @[MUL.scala 102:19]
  wire  m_2168_io_s; // @[MUL.scala 102:19]
  wire  m_2168_io_cout; // @[MUL.scala 102:19]
  wire  m_2169_io_x1; // @[MUL.scala 102:19]
  wire  m_2169_io_x2; // @[MUL.scala 102:19]
  wire  m_2169_io_x3; // @[MUL.scala 102:19]
  wire  m_2169_io_s; // @[MUL.scala 102:19]
  wire  m_2169_io_cout; // @[MUL.scala 102:19]
  wire  m_2170_io_x1; // @[MUL.scala 102:19]
  wire  m_2170_io_x2; // @[MUL.scala 102:19]
  wire  m_2170_io_x3; // @[MUL.scala 102:19]
  wire  m_2170_io_s; // @[MUL.scala 102:19]
  wire  m_2170_io_cout; // @[MUL.scala 102:19]
  wire  m_2171_io_x1; // @[MUL.scala 102:19]
  wire  m_2171_io_x2; // @[MUL.scala 102:19]
  wire  m_2171_io_x3; // @[MUL.scala 102:19]
  wire  m_2171_io_s; // @[MUL.scala 102:19]
  wire  m_2171_io_cout; // @[MUL.scala 102:19]
  wire  m_2172_io_x1; // @[MUL.scala 102:19]
  wire  m_2172_io_x2; // @[MUL.scala 102:19]
  wire  m_2172_io_x3; // @[MUL.scala 102:19]
  wire  m_2172_io_s; // @[MUL.scala 102:19]
  wire  m_2172_io_cout; // @[MUL.scala 102:19]
  wire  m_2173_io_x1; // @[MUL.scala 102:19]
  wire  m_2173_io_x2; // @[MUL.scala 102:19]
  wire  m_2173_io_x3; // @[MUL.scala 102:19]
  wire  m_2173_io_s; // @[MUL.scala 102:19]
  wire  m_2173_io_cout; // @[MUL.scala 102:19]
  wire  m_2174_io_x1; // @[MUL.scala 102:19]
  wire  m_2174_io_x2; // @[MUL.scala 102:19]
  wire  m_2174_io_x3; // @[MUL.scala 102:19]
  wire  m_2174_io_s; // @[MUL.scala 102:19]
  wire  m_2174_io_cout; // @[MUL.scala 102:19]
  wire  m_2175_io_x1; // @[MUL.scala 102:19]
  wire  m_2175_io_x2; // @[MUL.scala 102:19]
  wire  m_2175_io_x3; // @[MUL.scala 102:19]
  wire  m_2175_io_s; // @[MUL.scala 102:19]
  wire  m_2175_io_cout; // @[MUL.scala 102:19]
  wire  m_2176_io_x1; // @[MUL.scala 102:19]
  wire  m_2176_io_x2; // @[MUL.scala 102:19]
  wire  m_2176_io_x3; // @[MUL.scala 102:19]
  wire  m_2176_io_s; // @[MUL.scala 102:19]
  wire  m_2176_io_cout; // @[MUL.scala 102:19]
  wire  m_2177_io_x1; // @[MUL.scala 102:19]
  wire  m_2177_io_x2; // @[MUL.scala 102:19]
  wire  m_2177_io_x3; // @[MUL.scala 102:19]
  wire  m_2177_io_s; // @[MUL.scala 102:19]
  wire  m_2177_io_cout; // @[MUL.scala 102:19]
  wire  m_2178_io_x1; // @[MUL.scala 102:19]
  wire  m_2178_io_x2; // @[MUL.scala 102:19]
  wire  m_2178_io_x3; // @[MUL.scala 102:19]
  wire  m_2178_io_s; // @[MUL.scala 102:19]
  wire  m_2178_io_cout; // @[MUL.scala 102:19]
  wire  m_2179_io_x1; // @[MUL.scala 102:19]
  wire  m_2179_io_x2; // @[MUL.scala 102:19]
  wire  m_2179_io_x3; // @[MUL.scala 102:19]
  wire  m_2179_io_s; // @[MUL.scala 102:19]
  wire  m_2179_io_cout; // @[MUL.scala 102:19]
  wire  m_2180_io_x1; // @[MUL.scala 102:19]
  wire  m_2180_io_x2; // @[MUL.scala 102:19]
  wire  m_2180_io_x3; // @[MUL.scala 102:19]
  wire  m_2180_io_s; // @[MUL.scala 102:19]
  wire  m_2180_io_cout; // @[MUL.scala 102:19]
  wire  m_2181_io_x1; // @[MUL.scala 102:19]
  wire  m_2181_io_x2; // @[MUL.scala 102:19]
  wire  m_2181_io_x3; // @[MUL.scala 102:19]
  wire  m_2181_io_s; // @[MUL.scala 102:19]
  wire  m_2181_io_cout; // @[MUL.scala 102:19]
  wire  m_2182_io_x1; // @[MUL.scala 102:19]
  wire  m_2182_io_x2; // @[MUL.scala 102:19]
  wire  m_2182_io_x3; // @[MUL.scala 102:19]
  wire  m_2182_io_s; // @[MUL.scala 102:19]
  wire  m_2182_io_cout; // @[MUL.scala 102:19]
  wire  m_2183_io_x1; // @[MUL.scala 102:19]
  wire  m_2183_io_x2; // @[MUL.scala 102:19]
  wire  m_2183_io_x3; // @[MUL.scala 102:19]
  wire  m_2183_io_s; // @[MUL.scala 102:19]
  wire  m_2183_io_cout; // @[MUL.scala 102:19]
  wire  m_2184_io_x1; // @[MUL.scala 102:19]
  wire  m_2184_io_x2; // @[MUL.scala 102:19]
  wire  m_2184_io_x3; // @[MUL.scala 102:19]
  wire  m_2184_io_s; // @[MUL.scala 102:19]
  wire  m_2184_io_cout; // @[MUL.scala 102:19]
  wire  m_2185_io_x1; // @[MUL.scala 102:19]
  wire  m_2185_io_x2; // @[MUL.scala 102:19]
  wire  m_2185_io_x3; // @[MUL.scala 102:19]
  wire  m_2185_io_s; // @[MUL.scala 102:19]
  wire  m_2185_io_cout; // @[MUL.scala 102:19]
  wire  m_2186_io_x1; // @[MUL.scala 102:19]
  wire  m_2186_io_x2; // @[MUL.scala 102:19]
  wire  m_2186_io_x3; // @[MUL.scala 102:19]
  wire  m_2186_io_s; // @[MUL.scala 102:19]
  wire  m_2186_io_cout; // @[MUL.scala 102:19]
  wire  m_2187_io_x1; // @[MUL.scala 102:19]
  wire  m_2187_io_x2; // @[MUL.scala 102:19]
  wire  m_2187_io_x3; // @[MUL.scala 102:19]
  wire  m_2187_io_s; // @[MUL.scala 102:19]
  wire  m_2187_io_cout; // @[MUL.scala 102:19]
  wire  m_2188_io_x1; // @[MUL.scala 102:19]
  wire  m_2188_io_x2; // @[MUL.scala 102:19]
  wire  m_2188_io_x3; // @[MUL.scala 102:19]
  wire  m_2188_io_s; // @[MUL.scala 102:19]
  wire  m_2188_io_cout; // @[MUL.scala 102:19]
  wire  m_2189_io_x1; // @[MUL.scala 102:19]
  wire  m_2189_io_x2; // @[MUL.scala 102:19]
  wire  m_2189_io_x3; // @[MUL.scala 102:19]
  wire  m_2189_io_s; // @[MUL.scala 102:19]
  wire  m_2189_io_cout; // @[MUL.scala 102:19]
  wire  m_2190_io_x1; // @[MUL.scala 102:19]
  wire  m_2190_io_x2; // @[MUL.scala 102:19]
  wire  m_2190_io_x3; // @[MUL.scala 102:19]
  wire  m_2190_io_s; // @[MUL.scala 102:19]
  wire  m_2190_io_cout; // @[MUL.scala 102:19]
  wire  m_2191_io_x1; // @[MUL.scala 102:19]
  wire  m_2191_io_x2; // @[MUL.scala 102:19]
  wire  m_2191_io_x3; // @[MUL.scala 102:19]
  wire  m_2191_io_s; // @[MUL.scala 102:19]
  wire  m_2191_io_cout; // @[MUL.scala 102:19]
  wire  m_2192_io_in_0; // @[MUL.scala 124:19]
  wire  m_2192_io_in_1; // @[MUL.scala 124:19]
  wire  m_2192_io_out_0; // @[MUL.scala 124:19]
  wire  m_2192_io_out_1; // @[MUL.scala 124:19]
  wire  m_2193_io_x1; // @[MUL.scala 102:19]
  wire  m_2193_io_x2; // @[MUL.scala 102:19]
  wire  m_2193_io_x3; // @[MUL.scala 102:19]
  wire  m_2193_io_s; // @[MUL.scala 102:19]
  wire  m_2193_io_cout; // @[MUL.scala 102:19]
  wire  m_2194_io_in_0; // @[MUL.scala 124:19]
  wire  m_2194_io_in_1; // @[MUL.scala 124:19]
  wire  m_2194_io_out_0; // @[MUL.scala 124:19]
  wire  m_2194_io_out_1; // @[MUL.scala 124:19]
  wire  m_2195_io_x1; // @[MUL.scala 102:19]
  wire  m_2195_io_x2; // @[MUL.scala 102:19]
  wire  m_2195_io_x3; // @[MUL.scala 102:19]
  wire  m_2195_io_s; // @[MUL.scala 102:19]
  wire  m_2195_io_cout; // @[MUL.scala 102:19]
  wire  m_2196_io_in_0; // @[MUL.scala 124:19]
  wire  m_2196_io_in_1; // @[MUL.scala 124:19]
  wire  m_2196_io_out_0; // @[MUL.scala 124:19]
  wire  m_2196_io_out_1; // @[MUL.scala 124:19]
  wire  m_2197_io_x1; // @[MUL.scala 102:19]
  wire  m_2197_io_x2; // @[MUL.scala 102:19]
  wire  m_2197_io_x3; // @[MUL.scala 102:19]
  wire  m_2197_io_s; // @[MUL.scala 102:19]
  wire  m_2197_io_cout; // @[MUL.scala 102:19]
  wire  m_2198_io_in_0; // @[MUL.scala 124:19]
  wire  m_2198_io_in_1; // @[MUL.scala 124:19]
  wire  m_2198_io_out_0; // @[MUL.scala 124:19]
  wire  m_2198_io_out_1; // @[MUL.scala 124:19]
  wire  m_2199_io_x1; // @[MUL.scala 102:19]
  wire  m_2199_io_x2; // @[MUL.scala 102:19]
  wire  m_2199_io_x3; // @[MUL.scala 102:19]
  wire  m_2199_io_s; // @[MUL.scala 102:19]
  wire  m_2199_io_cout; // @[MUL.scala 102:19]
  wire  m_2200_io_in_0; // @[MUL.scala 124:19]
  wire  m_2200_io_in_1; // @[MUL.scala 124:19]
  wire  m_2200_io_out_0; // @[MUL.scala 124:19]
  wire  m_2200_io_out_1; // @[MUL.scala 124:19]
  wire  m_2201_io_x1; // @[MUL.scala 102:19]
  wire  m_2201_io_x2; // @[MUL.scala 102:19]
  wire  m_2201_io_x3; // @[MUL.scala 102:19]
  wire  m_2201_io_s; // @[MUL.scala 102:19]
  wire  m_2201_io_cout; // @[MUL.scala 102:19]
  wire  m_2202_io_in_0; // @[MUL.scala 124:19]
  wire  m_2202_io_in_1; // @[MUL.scala 124:19]
  wire  m_2202_io_out_0; // @[MUL.scala 124:19]
  wire  m_2202_io_out_1; // @[MUL.scala 124:19]
  wire  m_2203_io_x1; // @[MUL.scala 102:19]
  wire  m_2203_io_x2; // @[MUL.scala 102:19]
  wire  m_2203_io_x3; // @[MUL.scala 102:19]
  wire  m_2203_io_s; // @[MUL.scala 102:19]
  wire  m_2203_io_cout; // @[MUL.scala 102:19]
  wire  m_2204_io_in_0; // @[MUL.scala 124:19]
  wire  m_2204_io_in_1; // @[MUL.scala 124:19]
  wire  m_2204_io_out_0; // @[MUL.scala 124:19]
  wire  m_2204_io_out_1; // @[MUL.scala 124:19]
  wire  m_2205_io_x1; // @[MUL.scala 102:19]
  wire  m_2205_io_x2; // @[MUL.scala 102:19]
  wire  m_2205_io_x3; // @[MUL.scala 102:19]
  wire  m_2205_io_s; // @[MUL.scala 102:19]
  wire  m_2205_io_cout; // @[MUL.scala 102:19]
  wire  m_2206_io_in_0; // @[MUL.scala 124:19]
  wire  m_2206_io_in_1; // @[MUL.scala 124:19]
  wire  m_2206_io_out_0; // @[MUL.scala 124:19]
  wire  m_2206_io_out_1; // @[MUL.scala 124:19]
  wire  m_2207_io_x1; // @[MUL.scala 102:19]
  wire  m_2207_io_x2; // @[MUL.scala 102:19]
  wire  m_2207_io_x3; // @[MUL.scala 102:19]
  wire  m_2207_io_s; // @[MUL.scala 102:19]
  wire  m_2207_io_cout; // @[MUL.scala 102:19]
  wire  m_2208_io_in_0; // @[MUL.scala 124:19]
  wire  m_2208_io_in_1; // @[MUL.scala 124:19]
  wire  m_2208_io_out_0; // @[MUL.scala 124:19]
  wire  m_2208_io_out_1; // @[MUL.scala 124:19]
  wire  m_2209_io_x1; // @[MUL.scala 102:19]
  wire  m_2209_io_x2; // @[MUL.scala 102:19]
  wire  m_2209_io_x3; // @[MUL.scala 102:19]
  wire  m_2209_io_s; // @[MUL.scala 102:19]
  wire  m_2209_io_cout; // @[MUL.scala 102:19]
  wire  m_2210_io_in_0; // @[MUL.scala 124:19]
  wire  m_2210_io_in_1; // @[MUL.scala 124:19]
  wire  m_2210_io_out_0; // @[MUL.scala 124:19]
  wire  m_2210_io_out_1; // @[MUL.scala 124:19]
  wire  m_2211_io_x1; // @[MUL.scala 102:19]
  wire  m_2211_io_x2; // @[MUL.scala 102:19]
  wire  m_2211_io_x3; // @[MUL.scala 102:19]
  wire  m_2211_io_s; // @[MUL.scala 102:19]
  wire  m_2211_io_cout; // @[MUL.scala 102:19]
  wire  m_2212_io_in_0; // @[MUL.scala 124:19]
  wire  m_2212_io_in_1; // @[MUL.scala 124:19]
  wire  m_2212_io_out_0; // @[MUL.scala 124:19]
  wire  m_2212_io_out_1; // @[MUL.scala 124:19]
  wire  m_2213_io_x1; // @[MUL.scala 102:19]
  wire  m_2213_io_x2; // @[MUL.scala 102:19]
  wire  m_2213_io_x3; // @[MUL.scala 102:19]
  wire  m_2213_io_s; // @[MUL.scala 102:19]
  wire  m_2213_io_cout; // @[MUL.scala 102:19]
  wire  m_2214_io_in_0; // @[MUL.scala 124:19]
  wire  m_2214_io_in_1; // @[MUL.scala 124:19]
  wire  m_2214_io_out_0; // @[MUL.scala 124:19]
  wire  m_2214_io_out_1; // @[MUL.scala 124:19]
  wire  m_2215_io_x1; // @[MUL.scala 102:19]
  wire  m_2215_io_x2; // @[MUL.scala 102:19]
  wire  m_2215_io_x3; // @[MUL.scala 102:19]
  wire  m_2215_io_s; // @[MUL.scala 102:19]
  wire  m_2215_io_cout; // @[MUL.scala 102:19]
  wire  m_2216_io_in_0; // @[MUL.scala 124:19]
  wire  m_2216_io_in_1; // @[MUL.scala 124:19]
  wire  m_2216_io_out_0; // @[MUL.scala 124:19]
  wire  m_2216_io_out_1; // @[MUL.scala 124:19]
  wire  m_2217_io_x1; // @[MUL.scala 102:19]
  wire  m_2217_io_x2; // @[MUL.scala 102:19]
  wire  m_2217_io_x3; // @[MUL.scala 102:19]
  wire  m_2217_io_s; // @[MUL.scala 102:19]
  wire  m_2217_io_cout; // @[MUL.scala 102:19]
  wire  m_2218_io_in_0; // @[MUL.scala 124:19]
  wire  m_2218_io_in_1; // @[MUL.scala 124:19]
  wire  m_2218_io_out_0; // @[MUL.scala 124:19]
  wire  m_2218_io_out_1; // @[MUL.scala 124:19]
  wire  m_2219_io_x1; // @[MUL.scala 102:19]
  wire  m_2219_io_x2; // @[MUL.scala 102:19]
  wire  m_2219_io_x3; // @[MUL.scala 102:19]
  wire  m_2219_io_s; // @[MUL.scala 102:19]
  wire  m_2219_io_cout; // @[MUL.scala 102:19]
  wire  m_2220_io_in_0; // @[MUL.scala 124:19]
  wire  m_2220_io_in_1; // @[MUL.scala 124:19]
  wire  m_2220_io_out_0; // @[MUL.scala 124:19]
  wire  m_2220_io_out_1; // @[MUL.scala 124:19]
  wire  m_2221_io_x1; // @[MUL.scala 102:19]
  wire  m_2221_io_x2; // @[MUL.scala 102:19]
  wire  m_2221_io_x3; // @[MUL.scala 102:19]
  wire  m_2221_io_s; // @[MUL.scala 102:19]
  wire  m_2221_io_cout; // @[MUL.scala 102:19]
  wire  m_2222_io_in_0; // @[MUL.scala 124:19]
  wire  m_2222_io_in_1; // @[MUL.scala 124:19]
  wire  m_2222_io_out_0; // @[MUL.scala 124:19]
  wire  m_2222_io_out_1; // @[MUL.scala 124:19]
  wire  m_2223_io_x1; // @[MUL.scala 102:19]
  wire  m_2223_io_x2; // @[MUL.scala 102:19]
  wire  m_2223_io_x3; // @[MUL.scala 102:19]
  wire  m_2223_io_s; // @[MUL.scala 102:19]
  wire  m_2223_io_cout; // @[MUL.scala 102:19]
  wire  m_2224_io_in_0; // @[MUL.scala 124:19]
  wire  m_2224_io_in_1; // @[MUL.scala 124:19]
  wire  m_2224_io_out_0; // @[MUL.scala 124:19]
  wire  m_2224_io_out_1; // @[MUL.scala 124:19]
  wire  m_2225_io_x1; // @[MUL.scala 102:19]
  wire  m_2225_io_x2; // @[MUL.scala 102:19]
  wire  m_2225_io_x3; // @[MUL.scala 102:19]
  wire  m_2225_io_s; // @[MUL.scala 102:19]
  wire  m_2225_io_cout; // @[MUL.scala 102:19]
  wire  m_2226_io_in_0; // @[MUL.scala 124:19]
  wire  m_2226_io_in_1; // @[MUL.scala 124:19]
  wire  m_2226_io_out_0; // @[MUL.scala 124:19]
  wire  m_2226_io_out_1; // @[MUL.scala 124:19]
  wire  m_2227_io_x1; // @[MUL.scala 102:19]
  wire  m_2227_io_x2; // @[MUL.scala 102:19]
  wire  m_2227_io_x3; // @[MUL.scala 102:19]
  wire  m_2227_io_s; // @[MUL.scala 102:19]
  wire  m_2227_io_cout; // @[MUL.scala 102:19]
  wire  m_2228_io_in_0; // @[MUL.scala 124:19]
  wire  m_2228_io_in_1; // @[MUL.scala 124:19]
  wire  m_2228_io_out_0; // @[MUL.scala 124:19]
  wire  m_2228_io_out_1; // @[MUL.scala 124:19]
  wire  m_2229_io_x1; // @[MUL.scala 102:19]
  wire  m_2229_io_x2; // @[MUL.scala 102:19]
  wire  m_2229_io_x3; // @[MUL.scala 102:19]
  wire  m_2229_io_s; // @[MUL.scala 102:19]
  wire  m_2229_io_cout; // @[MUL.scala 102:19]
  wire  m_2230_io_in_0; // @[MUL.scala 124:19]
  wire  m_2230_io_in_1; // @[MUL.scala 124:19]
  wire  m_2230_io_out_0; // @[MUL.scala 124:19]
  wire  m_2230_io_out_1; // @[MUL.scala 124:19]
  wire  m_2231_io_x1; // @[MUL.scala 102:19]
  wire  m_2231_io_x2; // @[MUL.scala 102:19]
  wire  m_2231_io_x3; // @[MUL.scala 102:19]
  wire  m_2231_io_s; // @[MUL.scala 102:19]
  wire  m_2231_io_cout; // @[MUL.scala 102:19]
  wire  m_2232_io_in_0; // @[MUL.scala 124:19]
  wire  m_2232_io_in_1; // @[MUL.scala 124:19]
  wire  m_2232_io_out_0; // @[MUL.scala 124:19]
  wire  m_2232_io_out_1; // @[MUL.scala 124:19]
  wire  m_2233_io_x1; // @[MUL.scala 102:19]
  wire  m_2233_io_x2; // @[MUL.scala 102:19]
  wire  m_2233_io_x3; // @[MUL.scala 102:19]
  wire  m_2233_io_s; // @[MUL.scala 102:19]
  wire  m_2233_io_cout; // @[MUL.scala 102:19]
  wire  m_2234_io_x1; // @[MUL.scala 102:19]
  wire  m_2234_io_x2; // @[MUL.scala 102:19]
  wire  m_2234_io_x3; // @[MUL.scala 102:19]
  wire  m_2234_io_s; // @[MUL.scala 102:19]
  wire  m_2234_io_cout; // @[MUL.scala 102:19]
  wire  m_2235_io_x1; // @[MUL.scala 102:19]
  wire  m_2235_io_x2; // @[MUL.scala 102:19]
  wire  m_2235_io_x3; // @[MUL.scala 102:19]
  wire  m_2235_io_s; // @[MUL.scala 102:19]
  wire  m_2235_io_cout; // @[MUL.scala 102:19]
  wire  m_2236_io_x1; // @[MUL.scala 102:19]
  wire  m_2236_io_x2; // @[MUL.scala 102:19]
  wire  m_2236_io_x3; // @[MUL.scala 102:19]
  wire  m_2236_io_s; // @[MUL.scala 102:19]
  wire  m_2236_io_cout; // @[MUL.scala 102:19]
  wire  m_2237_io_x1; // @[MUL.scala 102:19]
  wire  m_2237_io_x2; // @[MUL.scala 102:19]
  wire  m_2237_io_x3; // @[MUL.scala 102:19]
  wire  m_2237_io_s; // @[MUL.scala 102:19]
  wire  m_2237_io_cout; // @[MUL.scala 102:19]
  wire  m_2238_io_x1; // @[MUL.scala 102:19]
  wire  m_2238_io_x2; // @[MUL.scala 102:19]
  wire  m_2238_io_x3; // @[MUL.scala 102:19]
  wire  m_2238_io_s; // @[MUL.scala 102:19]
  wire  m_2238_io_cout; // @[MUL.scala 102:19]
  wire  m_2239_io_x1; // @[MUL.scala 102:19]
  wire  m_2239_io_x2; // @[MUL.scala 102:19]
  wire  m_2239_io_x3; // @[MUL.scala 102:19]
  wire  m_2239_io_s; // @[MUL.scala 102:19]
  wire  m_2239_io_cout; // @[MUL.scala 102:19]
  wire  m_2240_io_x1; // @[MUL.scala 102:19]
  wire  m_2240_io_x2; // @[MUL.scala 102:19]
  wire  m_2240_io_x3; // @[MUL.scala 102:19]
  wire  m_2240_io_s; // @[MUL.scala 102:19]
  wire  m_2240_io_cout; // @[MUL.scala 102:19]
  wire  m_2241_io_x1; // @[MUL.scala 102:19]
  wire  m_2241_io_x2; // @[MUL.scala 102:19]
  wire  m_2241_io_x3; // @[MUL.scala 102:19]
  wire  m_2241_io_s; // @[MUL.scala 102:19]
  wire  m_2241_io_cout; // @[MUL.scala 102:19]
  wire  m_2242_io_x1; // @[MUL.scala 102:19]
  wire  m_2242_io_x2; // @[MUL.scala 102:19]
  wire  m_2242_io_x3; // @[MUL.scala 102:19]
  wire  m_2242_io_s; // @[MUL.scala 102:19]
  wire  m_2242_io_cout; // @[MUL.scala 102:19]
  wire  m_2243_io_x1; // @[MUL.scala 102:19]
  wire  m_2243_io_x2; // @[MUL.scala 102:19]
  wire  m_2243_io_x3; // @[MUL.scala 102:19]
  wire  m_2243_io_s; // @[MUL.scala 102:19]
  wire  m_2243_io_cout; // @[MUL.scala 102:19]
  wire  m_2244_io_x1; // @[MUL.scala 102:19]
  wire  m_2244_io_x2; // @[MUL.scala 102:19]
  wire  m_2244_io_x3; // @[MUL.scala 102:19]
  wire  m_2244_io_s; // @[MUL.scala 102:19]
  wire  m_2244_io_cout; // @[MUL.scala 102:19]
  wire  m_2245_io_x1; // @[MUL.scala 102:19]
  wire  m_2245_io_x2; // @[MUL.scala 102:19]
  wire  m_2245_io_x3; // @[MUL.scala 102:19]
  wire  m_2245_io_s; // @[MUL.scala 102:19]
  wire  m_2245_io_cout; // @[MUL.scala 102:19]
  wire  m_2246_io_x1; // @[MUL.scala 102:19]
  wire  m_2246_io_x2; // @[MUL.scala 102:19]
  wire  m_2246_io_x3; // @[MUL.scala 102:19]
  wire  m_2246_io_s; // @[MUL.scala 102:19]
  wire  m_2246_io_cout; // @[MUL.scala 102:19]
  wire  m_2247_io_x1; // @[MUL.scala 102:19]
  wire  m_2247_io_x2; // @[MUL.scala 102:19]
  wire  m_2247_io_x3; // @[MUL.scala 102:19]
  wire  m_2247_io_s; // @[MUL.scala 102:19]
  wire  m_2247_io_cout; // @[MUL.scala 102:19]
  wire  m_2248_io_x1; // @[MUL.scala 102:19]
  wire  m_2248_io_x2; // @[MUL.scala 102:19]
  wire  m_2248_io_x3; // @[MUL.scala 102:19]
  wire  m_2248_io_s; // @[MUL.scala 102:19]
  wire  m_2248_io_cout; // @[MUL.scala 102:19]
  wire  m_2249_io_x1; // @[MUL.scala 102:19]
  wire  m_2249_io_x2; // @[MUL.scala 102:19]
  wire  m_2249_io_x3; // @[MUL.scala 102:19]
  wire  m_2249_io_s; // @[MUL.scala 102:19]
  wire  m_2249_io_cout; // @[MUL.scala 102:19]
  wire  m_2250_io_x1; // @[MUL.scala 102:19]
  wire  m_2250_io_x2; // @[MUL.scala 102:19]
  wire  m_2250_io_x3; // @[MUL.scala 102:19]
  wire  m_2250_io_s; // @[MUL.scala 102:19]
  wire  m_2250_io_cout; // @[MUL.scala 102:19]
  wire  m_2251_io_x1; // @[MUL.scala 102:19]
  wire  m_2251_io_x2; // @[MUL.scala 102:19]
  wire  m_2251_io_x3; // @[MUL.scala 102:19]
  wire  m_2251_io_s; // @[MUL.scala 102:19]
  wire  m_2251_io_cout; // @[MUL.scala 102:19]
  wire  m_2252_io_x1; // @[MUL.scala 102:19]
  wire  m_2252_io_x2; // @[MUL.scala 102:19]
  wire  m_2252_io_x3; // @[MUL.scala 102:19]
  wire  m_2252_io_s; // @[MUL.scala 102:19]
  wire  m_2252_io_cout; // @[MUL.scala 102:19]
  wire  m_2253_io_x1; // @[MUL.scala 102:19]
  wire  m_2253_io_x2; // @[MUL.scala 102:19]
  wire  m_2253_io_x3; // @[MUL.scala 102:19]
  wire  m_2253_io_s; // @[MUL.scala 102:19]
  wire  m_2253_io_cout; // @[MUL.scala 102:19]
  wire  m_2254_io_x1; // @[MUL.scala 102:19]
  wire  m_2254_io_x2; // @[MUL.scala 102:19]
  wire  m_2254_io_x3; // @[MUL.scala 102:19]
  wire  m_2254_io_s; // @[MUL.scala 102:19]
  wire  m_2254_io_cout; // @[MUL.scala 102:19]
  wire  m_2255_io_x1; // @[MUL.scala 102:19]
  wire  m_2255_io_x2; // @[MUL.scala 102:19]
  wire  m_2255_io_x3; // @[MUL.scala 102:19]
  wire  m_2255_io_s; // @[MUL.scala 102:19]
  wire  m_2255_io_cout; // @[MUL.scala 102:19]
  wire  m_2256_io_x1; // @[MUL.scala 102:19]
  wire  m_2256_io_x2; // @[MUL.scala 102:19]
  wire  m_2256_io_x3; // @[MUL.scala 102:19]
  wire  m_2256_io_s; // @[MUL.scala 102:19]
  wire  m_2256_io_cout; // @[MUL.scala 102:19]
  wire  m_2257_io_x1; // @[MUL.scala 102:19]
  wire  m_2257_io_x2; // @[MUL.scala 102:19]
  wire  m_2257_io_x3; // @[MUL.scala 102:19]
  wire  m_2257_io_s; // @[MUL.scala 102:19]
  wire  m_2257_io_cout; // @[MUL.scala 102:19]
  wire  m_2258_io_x1; // @[MUL.scala 102:19]
  wire  m_2258_io_x2; // @[MUL.scala 102:19]
  wire  m_2258_io_x3; // @[MUL.scala 102:19]
  wire  m_2258_io_s; // @[MUL.scala 102:19]
  wire  m_2258_io_cout; // @[MUL.scala 102:19]
  wire  m_2259_io_x1; // @[MUL.scala 102:19]
  wire  m_2259_io_x2; // @[MUL.scala 102:19]
  wire  m_2259_io_x3; // @[MUL.scala 102:19]
  wire  m_2259_io_s; // @[MUL.scala 102:19]
  wire  m_2259_io_cout; // @[MUL.scala 102:19]
  wire  m_2260_io_x1; // @[MUL.scala 102:19]
  wire  m_2260_io_x2; // @[MUL.scala 102:19]
  wire  m_2260_io_x3; // @[MUL.scala 102:19]
  wire  m_2260_io_s; // @[MUL.scala 102:19]
  wire  m_2260_io_cout; // @[MUL.scala 102:19]
  wire  m_2261_io_x1; // @[MUL.scala 102:19]
  wire  m_2261_io_x2; // @[MUL.scala 102:19]
  wire  m_2261_io_x3; // @[MUL.scala 102:19]
  wire  m_2261_io_s; // @[MUL.scala 102:19]
  wire  m_2261_io_cout; // @[MUL.scala 102:19]
  wire  m_2262_io_x1; // @[MUL.scala 102:19]
  wire  m_2262_io_x2; // @[MUL.scala 102:19]
  wire  m_2262_io_x3; // @[MUL.scala 102:19]
  wire  m_2262_io_s; // @[MUL.scala 102:19]
  wire  m_2262_io_cout; // @[MUL.scala 102:19]
  wire  m_2263_io_in_0; // @[MUL.scala 124:19]
  wire  m_2263_io_in_1; // @[MUL.scala 124:19]
  wire  m_2263_io_out_0; // @[MUL.scala 124:19]
  wire  m_2263_io_out_1; // @[MUL.scala 124:19]
  wire  m_2264_io_in_0; // @[MUL.scala 124:19]
  wire  m_2264_io_in_1; // @[MUL.scala 124:19]
  wire  m_2264_io_out_0; // @[MUL.scala 124:19]
  wire  m_2264_io_out_1; // @[MUL.scala 124:19]
  wire  m_2265_io_in_0; // @[MUL.scala 124:19]
  wire  m_2265_io_in_1; // @[MUL.scala 124:19]
  wire  m_2265_io_out_0; // @[MUL.scala 124:19]
  wire  m_2265_io_out_1; // @[MUL.scala 124:19]
  wire  m_2266_io_in_0; // @[MUL.scala 124:19]
  wire  m_2266_io_in_1; // @[MUL.scala 124:19]
  wire  m_2266_io_out_0; // @[MUL.scala 124:19]
  wire  m_2266_io_out_1; // @[MUL.scala 124:19]
  wire  m_2267_io_in_0; // @[MUL.scala 124:19]
  wire  m_2267_io_in_1; // @[MUL.scala 124:19]
  wire  m_2267_io_out_0; // @[MUL.scala 124:19]
  wire  m_2267_io_out_1; // @[MUL.scala 124:19]
  wire  m_2268_io_in_0; // @[MUL.scala 124:19]
  wire  m_2268_io_in_1; // @[MUL.scala 124:19]
  wire  m_2268_io_out_0; // @[MUL.scala 124:19]
  wire  m_2268_io_out_1; // @[MUL.scala 124:19]
  wire  m_2269_io_in_0; // @[MUL.scala 124:19]
  wire  m_2269_io_in_1; // @[MUL.scala 124:19]
  wire  m_2269_io_out_0; // @[MUL.scala 124:19]
  wire  m_2269_io_out_1; // @[MUL.scala 124:19]
  wire  m_2270_io_in_0; // @[MUL.scala 124:19]
  wire  m_2270_io_in_1; // @[MUL.scala 124:19]
  wire  m_2270_io_out_0; // @[MUL.scala 124:19]
  wire  m_2270_io_out_1; // @[MUL.scala 124:19]
  wire  m_2271_io_in_0; // @[MUL.scala 124:19]
  wire  m_2271_io_in_1; // @[MUL.scala 124:19]
  wire  m_2271_io_out_0; // @[MUL.scala 124:19]
  wire  m_2271_io_out_1; // @[MUL.scala 124:19]
  wire  m_2272_io_in_0; // @[MUL.scala 124:19]
  wire  m_2272_io_in_1; // @[MUL.scala 124:19]
  wire  m_2272_io_out_0; // @[MUL.scala 124:19]
  wire  m_2272_io_out_1; // @[MUL.scala 124:19]
  wire  m_2273_io_in_0; // @[MUL.scala 124:19]
  wire  m_2273_io_in_1; // @[MUL.scala 124:19]
  wire  m_2273_io_out_0; // @[MUL.scala 124:19]
  wire  m_2273_io_out_1; // @[MUL.scala 124:19]
  wire  m_2274_io_in_0; // @[MUL.scala 124:19]
  wire  m_2274_io_in_1; // @[MUL.scala 124:19]
  wire  m_2274_io_out_0; // @[MUL.scala 124:19]
  wire  m_2274_io_out_1; // @[MUL.scala 124:19]
  wire  m_2275_io_in_0; // @[MUL.scala 124:19]
  wire  m_2275_io_in_1; // @[MUL.scala 124:19]
  wire  m_2275_io_out_0; // @[MUL.scala 124:19]
  wire  m_2275_io_out_1; // @[MUL.scala 124:19]
  wire  m_2276_io_in_0; // @[MUL.scala 124:19]
  wire  m_2276_io_in_1; // @[MUL.scala 124:19]
  wire  m_2276_io_out_0; // @[MUL.scala 124:19]
  wire  m_2276_io_out_1; // @[MUL.scala 124:19]
  wire  m_2277_io_in_0; // @[MUL.scala 124:19]
  wire  m_2277_io_in_1; // @[MUL.scala 124:19]
  wire  m_2277_io_out_0; // @[MUL.scala 124:19]
  wire  m_2277_io_out_1; // @[MUL.scala 124:19]
  wire  m_2278_io_in_0; // @[MUL.scala 124:19]
  wire  m_2278_io_in_1; // @[MUL.scala 124:19]
  wire  m_2278_io_out_0; // @[MUL.scala 124:19]
  wire  m_2278_io_out_1; // @[MUL.scala 124:19]
  wire  m_2279_io_in_0; // @[MUL.scala 124:19]
  wire  m_2279_io_in_1; // @[MUL.scala 124:19]
  wire  m_2279_io_out_0; // @[MUL.scala 124:19]
  wire  m_2279_io_out_1; // @[MUL.scala 124:19]
  wire  m_2280_io_in_0; // @[MUL.scala 124:19]
  wire  m_2280_io_in_1; // @[MUL.scala 124:19]
  wire  m_2280_io_out_0; // @[MUL.scala 124:19]
  wire  m_2280_io_out_1; // @[MUL.scala 124:19]
  wire  m_2281_io_in_0; // @[MUL.scala 124:19]
  wire  m_2281_io_in_1; // @[MUL.scala 124:19]
  wire  m_2281_io_out_0; // @[MUL.scala 124:19]
  wire  m_2281_io_out_1; // @[MUL.scala 124:19]
  wire  m_2282_io_in_0; // @[MUL.scala 124:19]
  wire  m_2282_io_in_1; // @[MUL.scala 124:19]
  wire  m_2282_io_out_0; // @[MUL.scala 124:19]
  wire  m_2282_io_out_1; // @[MUL.scala 124:19]
  wire  m_2283_io_in_0; // @[MUL.scala 124:19]
  wire  m_2283_io_in_1; // @[MUL.scala 124:19]
  wire  m_2283_io_out_0; // @[MUL.scala 124:19]
  wire  m_2283_io_out_1; // @[MUL.scala 124:19]
  wire  m_2284_io_in_0; // @[MUL.scala 124:19]
  wire  m_2284_io_in_1; // @[MUL.scala 124:19]
  wire  m_2284_io_out_0; // @[MUL.scala 124:19]
  wire  m_2284_io_out_1; // @[MUL.scala 124:19]
  wire  m_2285_io_in_0; // @[MUL.scala 124:19]
  wire  m_2285_io_in_1; // @[MUL.scala 124:19]
  wire  m_2285_io_out_0; // @[MUL.scala 124:19]
  wire  m_2285_io_out_1; // @[MUL.scala 124:19]
  wire  m_2286_io_in_0; // @[MUL.scala 124:19]
  wire  m_2286_io_in_1; // @[MUL.scala 124:19]
  wire  m_2286_io_out_0; // @[MUL.scala 124:19]
  wire  m_2286_io_out_1; // @[MUL.scala 124:19]
  wire  m_2287_io_in_0; // @[MUL.scala 124:19]
  wire  m_2287_io_in_1; // @[MUL.scala 124:19]
  wire  m_2287_io_out_0; // @[MUL.scala 124:19]
  wire  m_2287_io_out_1; // @[MUL.scala 124:19]
  wire  m_2288_io_in_0; // @[MUL.scala 124:19]
  wire  m_2288_io_in_1; // @[MUL.scala 124:19]
  wire  m_2288_io_out_0; // @[MUL.scala 124:19]
  wire  m_2288_io_out_1; // @[MUL.scala 124:19]
  wire  m_2289_io_in_0; // @[MUL.scala 124:19]
  wire  m_2289_io_in_1; // @[MUL.scala 124:19]
  wire  m_2289_io_out_0; // @[MUL.scala 124:19]
  wire  m_2289_io_out_1; // @[MUL.scala 124:19]
  wire  m_2290_io_in_0; // @[MUL.scala 124:19]
  wire  m_2290_io_in_1; // @[MUL.scala 124:19]
  wire  m_2290_io_out_0; // @[MUL.scala 124:19]
  wire  m_2290_io_out_1; // @[MUL.scala 124:19]
  wire  m_2291_io_in_0; // @[MUL.scala 124:19]
  wire  m_2291_io_in_1; // @[MUL.scala 124:19]
  wire  m_2291_io_out_0; // @[MUL.scala 124:19]
  wire  m_2291_io_out_1; // @[MUL.scala 124:19]
  wire  m_2292_io_in_0; // @[MUL.scala 124:19]
  wire  m_2292_io_in_1; // @[MUL.scala 124:19]
  wire  m_2292_io_out_0; // @[MUL.scala 124:19]
  wire  m_2292_io_out_1; // @[MUL.scala 124:19]
  wire  m_2293_io_in_0; // @[MUL.scala 124:19]
  wire  m_2293_io_in_1; // @[MUL.scala 124:19]
  wire  m_2293_io_out_0; // @[MUL.scala 124:19]
  wire  m_2293_io_out_1; // @[MUL.scala 124:19]
  wire  m_2294_io_in_0; // @[MUL.scala 124:19]
  wire  m_2294_io_in_1; // @[MUL.scala 124:19]
  wire  m_2294_io_out_0; // @[MUL.scala 124:19]
  wire  m_2294_io_out_1; // @[MUL.scala 124:19]
  wire  m_2295_io_in_0; // @[MUL.scala 124:19]
  wire  m_2295_io_in_1; // @[MUL.scala 124:19]
  wire  m_2295_io_out_0; // @[MUL.scala 124:19]
  wire  m_2295_io_out_1; // @[MUL.scala 124:19]
  wire  m_2296_io_in_0; // @[MUL.scala 124:19]
  wire  m_2296_io_in_1; // @[MUL.scala 124:19]
  wire  m_2296_io_out_0; // @[MUL.scala 124:19]
  wire  m_2296_io_out_1; // @[MUL.scala 124:19]
  wire  m_2297_io_in_0; // @[MUL.scala 124:19]
  wire  m_2297_io_in_1; // @[MUL.scala 124:19]
  wire  m_2297_io_out_0; // @[MUL.scala 124:19]
  wire  m_2297_io_out_1; // @[MUL.scala 124:19]
  wire  m_2298_io_in_0; // @[MUL.scala 124:19]
  wire  m_2298_io_in_1; // @[MUL.scala 124:19]
  wire  m_2298_io_out_0; // @[MUL.scala 124:19]
  wire  m_2298_io_out_1; // @[MUL.scala 124:19]
  wire  m_2299_io_in_0; // @[MUL.scala 124:19]
  wire  m_2299_io_in_1; // @[MUL.scala 124:19]
  wire  m_2299_io_out_0; // @[MUL.scala 124:19]
  wire  m_2299_io_out_1; // @[MUL.scala 124:19]
  wire  m_2300_io_in_0; // @[MUL.scala 124:19]
  wire  m_2300_io_in_1; // @[MUL.scala 124:19]
  wire  m_2300_io_out_0; // @[MUL.scala 124:19]
  wire  m_2300_io_out_1; // @[MUL.scala 124:19]
  wire  m_2301_io_in_0; // @[MUL.scala 124:19]
  wire  m_2301_io_in_1; // @[MUL.scala 124:19]
  wire  m_2301_io_out_0; // @[MUL.scala 124:19]
  wire  m_2301_io_out_1; // @[MUL.scala 124:19]
  wire  m_2302_io_in_0; // @[MUL.scala 124:19]
  wire  m_2302_io_in_1; // @[MUL.scala 124:19]
  wire  m_2302_io_out_0; // @[MUL.scala 124:19]
  wire  m_2302_io_out_1; // @[MUL.scala 124:19]
  wire  m_2303_io_in_0; // @[MUL.scala 124:19]
  wire  m_2303_io_in_1; // @[MUL.scala 124:19]
  wire  m_2303_io_out_0; // @[MUL.scala 124:19]
  wire  m_2303_io_out_1; // @[MUL.scala 124:19]
  wire  m_2304_io_in_0; // @[MUL.scala 124:19]
  wire  m_2304_io_in_1; // @[MUL.scala 124:19]
  wire  m_2304_io_out_0; // @[MUL.scala 124:19]
  wire  m_2304_io_out_1; // @[MUL.scala 124:19]
  wire  m_2305_io_in_0; // @[MUL.scala 124:19]
  wire  m_2305_io_in_1; // @[MUL.scala 124:19]
  wire  m_2305_io_out_0; // @[MUL.scala 124:19]
  wire  m_2305_io_out_1; // @[MUL.scala 124:19]
  wire  m_2306_io_in_0; // @[MUL.scala 124:19]
  wire  m_2306_io_in_1; // @[MUL.scala 124:19]
  wire  m_2306_io_out_0; // @[MUL.scala 124:19]
  wire  m_2306_io_out_1; // @[MUL.scala 124:19]
  wire  m_2307_io_in_0; // @[MUL.scala 124:19]
  wire  m_2307_io_in_1; // @[MUL.scala 124:19]
  wire  m_2307_io_out_0; // @[MUL.scala 124:19]
  wire  m_2307_io_out_1; // @[MUL.scala 124:19]
  wire  m_2308_io_in_0; // @[MUL.scala 124:19]
  wire  m_2308_io_in_1; // @[MUL.scala 124:19]
  wire  m_2308_io_out_0; // @[MUL.scala 124:19]
  wire  m_2308_io_out_1; // @[MUL.scala 124:19]
  wire  m_2309_io_in_0; // @[MUL.scala 124:19]
  wire  m_2309_io_in_1; // @[MUL.scala 124:19]
  wire  m_2309_io_out_0; // @[MUL.scala 124:19]
  wire  m_2309_io_out_1; // @[MUL.scala 124:19]
  wire  m_2310_io_in_0; // @[MUL.scala 124:19]
  wire  m_2310_io_in_1; // @[MUL.scala 124:19]
  wire  m_2310_io_out_0; // @[MUL.scala 124:19]
  wire  m_2310_io_out_1; // @[MUL.scala 124:19]
  wire  m_2311_io_in_0; // @[MUL.scala 124:19]
  wire  m_2311_io_in_1; // @[MUL.scala 124:19]
  wire  m_2311_io_out_0; // @[MUL.scala 124:19]
  wire  m_2311_io_out_1; // @[MUL.scala 124:19]
  wire  m_2312_io_in_0; // @[MUL.scala 124:19]
  wire  m_2312_io_in_1; // @[MUL.scala 124:19]
  wire  m_2312_io_out_0; // @[MUL.scala 124:19]
  wire  m_2312_io_out_1; // @[MUL.scala 124:19]
  wire  m_2313_io_in_0; // @[MUL.scala 124:19]
  wire  m_2313_io_in_1; // @[MUL.scala 124:19]
  wire  m_2313_io_out_0; // @[MUL.scala 124:19]
  wire  m_2313_io_out_1; // @[MUL.scala 124:19]
  wire  m_2314_io_in_0; // @[MUL.scala 124:19]
  wire  m_2314_io_in_1; // @[MUL.scala 124:19]
  wire  m_2314_io_out_0; // @[MUL.scala 124:19]
  wire  m_2314_io_out_1; // @[MUL.scala 124:19]
  wire  m_2315_io_in_0; // @[MUL.scala 124:19]
  wire  m_2315_io_in_1; // @[MUL.scala 124:19]
  wire  m_2315_io_out_0; // @[MUL.scala 124:19]
  wire  m_2315_io_out_1; // @[MUL.scala 124:19]
  wire  m_2316_io_in_0; // @[MUL.scala 124:19]
  wire  m_2316_io_in_1; // @[MUL.scala 124:19]
  wire  m_2316_io_out_0; // @[MUL.scala 124:19]
  wire  m_2316_io_out_1; // @[MUL.scala 124:19]
  wire  m_2317_io_in_0; // @[MUL.scala 124:19]
  wire  m_2317_io_in_1; // @[MUL.scala 124:19]
  wire  m_2317_io_out_0; // @[MUL.scala 124:19]
  wire  m_2317_io_out_1; // @[MUL.scala 124:19]
  wire  m_2318_io_in_0; // @[MUL.scala 124:19]
  wire  m_2318_io_in_1; // @[MUL.scala 124:19]
  wire  m_2318_io_out_0; // @[MUL.scala 124:19]
  wire  m_2318_io_out_1; // @[MUL.scala 124:19]
  wire  m_2319_io_x1; // @[MUL.scala 102:19]
  wire  m_2319_io_x2; // @[MUL.scala 102:19]
  wire  m_2319_io_x3; // @[MUL.scala 102:19]
  wire  m_2319_io_s; // @[MUL.scala 102:19]
  wire  m_2319_io_cout; // @[MUL.scala 102:19]
  wire  m_2320_io_x1; // @[MUL.scala 102:19]
  wire  m_2320_io_x2; // @[MUL.scala 102:19]
  wire  m_2320_io_x3; // @[MUL.scala 102:19]
  wire  m_2320_io_s; // @[MUL.scala 102:19]
  wire  m_2320_io_cout; // @[MUL.scala 102:19]
  wire  m_2321_io_x1; // @[MUL.scala 102:19]
  wire  m_2321_io_x2; // @[MUL.scala 102:19]
  wire  m_2321_io_x3; // @[MUL.scala 102:19]
  wire  m_2321_io_s; // @[MUL.scala 102:19]
  wire  m_2321_io_cout; // @[MUL.scala 102:19]
  wire  m_2322_io_x1; // @[MUL.scala 102:19]
  wire  m_2322_io_x2; // @[MUL.scala 102:19]
  wire  m_2322_io_x3; // @[MUL.scala 102:19]
  wire  m_2322_io_s; // @[MUL.scala 102:19]
  wire  m_2322_io_cout; // @[MUL.scala 102:19]
  wire  m_2323_io_x1; // @[MUL.scala 102:19]
  wire  m_2323_io_x2; // @[MUL.scala 102:19]
  wire  m_2323_io_x3; // @[MUL.scala 102:19]
  wire  m_2323_io_s; // @[MUL.scala 102:19]
  wire  m_2323_io_cout; // @[MUL.scala 102:19]
  wire  m_2324_io_x1; // @[MUL.scala 102:19]
  wire  m_2324_io_x2; // @[MUL.scala 102:19]
  wire  m_2324_io_x3; // @[MUL.scala 102:19]
  wire  m_2324_io_s; // @[MUL.scala 102:19]
  wire  m_2324_io_cout; // @[MUL.scala 102:19]
  wire  m_2325_io_x1; // @[MUL.scala 102:19]
  wire  m_2325_io_x2; // @[MUL.scala 102:19]
  wire  m_2325_io_x3; // @[MUL.scala 102:19]
  wire  m_2325_io_s; // @[MUL.scala 102:19]
  wire  m_2325_io_cout; // @[MUL.scala 102:19]
  wire  m_2326_io_x1; // @[MUL.scala 102:19]
  wire  m_2326_io_x2; // @[MUL.scala 102:19]
  wire  m_2326_io_x3; // @[MUL.scala 102:19]
  wire  m_2326_io_s; // @[MUL.scala 102:19]
  wire  m_2326_io_cout; // @[MUL.scala 102:19]
  wire  m_2327_io_x1; // @[MUL.scala 102:19]
  wire  m_2327_io_x2; // @[MUL.scala 102:19]
  wire  m_2327_io_x3; // @[MUL.scala 102:19]
  wire  m_2327_io_s; // @[MUL.scala 102:19]
  wire  m_2327_io_cout; // @[MUL.scala 102:19]
  wire  m_2328_io_x1; // @[MUL.scala 102:19]
  wire  m_2328_io_x2; // @[MUL.scala 102:19]
  wire  m_2328_io_x3; // @[MUL.scala 102:19]
  wire  m_2328_io_s; // @[MUL.scala 102:19]
  wire  m_2328_io_cout; // @[MUL.scala 102:19]
  wire  m_2329_io_x1; // @[MUL.scala 102:19]
  wire  m_2329_io_x2; // @[MUL.scala 102:19]
  wire  m_2329_io_x3; // @[MUL.scala 102:19]
  wire  m_2329_io_s; // @[MUL.scala 102:19]
  wire  m_2329_io_cout; // @[MUL.scala 102:19]
  wire  m_2330_io_x1; // @[MUL.scala 102:19]
  wire  m_2330_io_x2; // @[MUL.scala 102:19]
  wire  m_2330_io_x3; // @[MUL.scala 102:19]
  wire  m_2330_io_s; // @[MUL.scala 102:19]
  wire  m_2330_io_cout; // @[MUL.scala 102:19]
  wire  m_2331_io_x1; // @[MUL.scala 102:19]
  wire  m_2331_io_x2; // @[MUL.scala 102:19]
  wire  m_2331_io_x3; // @[MUL.scala 102:19]
  wire  m_2331_io_s; // @[MUL.scala 102:19]
  wire  m_2331_io_cout; // @[MUL.scala 102:19]
  wire  m_2332_io_x1; // @[MUL.scala 102:19]
  wire  m_2332_io_x2; // @[MUL.scala 102:19]
  wire  m_2332_io_x3; // @[MUL.scala 102:19]
  wire  m_2332_io_s; // @[MUL.scala 102:19]
  wire  m_2332_io_cout; // @[MUL.scala 102:19]
  wire  m_2333_io_x1; // @[MUL.scala 102:19]
  wire  m_2333_io_x2; // @[MUL.scala 102:19]
  wire  m_2333_io_x3; // @[MUL.scala 102:19]
  wire  m_2333_io_s; // @[MUL.scala 102:19]
  wire  m_2333_io_cout; // @[MUL.scala 102:19]
  wire  m_2334_io_x1; // @[MUL.scala 102:19]
  wire  m_2334_io_x2; // @[MUL.scala 102:19]
  wire  m_2334_io_x3; // @[MUL.scala 102:19]
  wire  m_2334_io_s; // @[MUL.scala 102:19]
  wire  m_2334_io_cout; // @[MUL.scala 102:19]
  wire  m_2335_io_x1; // @[MUL.scala 102:19]
  wire  m_2335_io_x2; // @[MUL.scala 102:19]
  wire  m_2335_io_x3; // @[MUL.scala 102:19]
  wire  m_2335_io_s; // @[MUL.scala 102:19]
  wire  m_2335_io_cout; // @[MUL.scala 102:19]
  wire  m_2336_io_x1; // @[MUL.scala 102:19]
  wire  m_2336_io_x2; // @[MUL.scala 102:19]
  wire  m_2336_io_x3; // @[MUL.scala 102:19]
  wire  m_2336_io_s; // @[MUL.scala 102:19]
  wire  m_2336_io_cout; // @[MUL.scala 102:19]
  wire  m_2337_io_x1; // @[MUL.scala 102:19]
  wire  m_2337_io_x2; // @[MUL.scala 102:19]
  wire  m_2337_io_x3; // @[MUL.scala 102:19]
  wire  m_2337_io_s; // @[MUL.scala 102:19]
  wire  m_2337_io_cout; // @[MUL.scala 102:19]
  wire  m_2338_io_x1; // @[MUL.scala 102:19]
  wire  m_2338_io_x2; // @[MUL.scala 102:19]
  wire  m_2338_io_x3; // @[MUL.scala 102:19]
  wire  m_2338_io_s; // @[MUL.scala 102:19]
  wire  m_2338_io_cout; // @[MUL.scala 102:19]
  wire  m_2339_io_x1; // @[MUL.scala 102:19]
  wire  m_2339_io_x2; // @[MUL.scala 102:19]
  wire  m_2339_io_x3; // @[MUL.scala 102:19]
  wire  m_2339_io_s; // @[MUL.scala 102:19]
  wire  m_2339_io_cout; // @[MUL.scala 102:19]
  wire  m_2340_io_x1; // @[MUL.scala 102:19]
  wire  m_2340_io_x2; // @[MUL.scala 102:19]
  wire  m_2340_io_x3; // @[MUL.scala 102:19]
  wire  m_2340_io_s; // @[MUL.scala 102:19]
  wire  m_2340_io_cout; // @[MUL.scala 102:19]
  wire  m_2341_io_x1; // @[MUL.scala 102:19]
  wire  m_2341_io_x2; // @[MUL.scala 102:19]
  wire  m_2341_io_x3; // @[MUL.scala 102:19]
  wire  m_2341_io_s; // @[MUL.scala 102:19]
  wire  m_2341_io_cout; // @[MUL.scala 102:19]
  wire  m_2342_io_x1; // @[MUL.scala 102:19]
  wire  m_2342_io_x2; // @[MUL.scala 102:19]
  wire  m_2342_io_x3; // @[MUL.scala 102:19]
  wire  m_2342_io_s; // @[MUL.scala 102:19]
  wire  m_2342_io_cout; // @[MUL.scala 102:19]
  wire  m_2343_io_x1; // @[MUL.scala 102:19]
  wire  m_2343_io_x2; // @[MUL.scala 102:19]
  wire  m_2343_io_x3; // @[MUL.scala 102:19]
  wire  m_2343_io_s; // @[MUL.scala 102:19]
  wire  m_2343_io_cout; // @[MUL.scala 102:19]
  wire  m_2344_io_x1; // @[MUL.scala 102:19]
  wire  m_2344_io_x2; // @[MUL.scala 102:19]
  wire  m_2344_io_x3; // @[MUL.scala 102:19]
  wire  m_2344_io_s; // @[MUL.scala 102:19]
  wire  m_2344_io_cout; // @[MUL.scala 102:19]
  wire  m_2345_io_x1; // @[MUL.scala 102:19]
  wire  m_2345_io_x2; // @[MUL.scala 102:19]
  wire  m_2345_io_x3; // @[MUL.scala 102:19]
  wire  m_2345_io_s; // @[MUL.scala 102:19]
  wire  m_2345_io_cout; // @[MUL.scala 102:19]
  wire  m_2346_io_x1; // @[MUL.scala 102:19]
  wire  m_2346_io_x2; // @[MUL.scala 102:19]
  wire  m_2346_io_x3; // @[MUL.scala 102:19]
  wire  m_2346_io_s; // @[MUL.scala 102:19]
  wire  m_2346_io_cout; // @[MUL.scala 102:19]
  wire  m_2347_io_x1; // @[MUL.scala 102:19]
  wire  m_2347_io_x2; // @[MUL.scala 102:19]
  wire  m_2347_io_x3; // @[MUL.scala 102:19]
  wire  m_2347_io_s; // @[MUL.scala 102:19]
  wire  m_2347_io_cout; // @[MUL.scala 102:19]
  wire  m_2348_io_x1; // @[MUL.scala 102:19]
  wire  m_2348_io_x2; // @[MUL.scala 102:19]
  wire  m_2348_io_x3; // @[MUL.scala 102:19]
  wire  m_2348_io_s; // @[MUL.scala 102:19]
  wire  m_2348_io_cout; // @[MUL.scala 102:19]
  wire  m_2349_io_x1; // @[MUL.scala 102:19]
  wire  m_2349_io_x2; // @[MUL.scala 102:19]
  wire  m_2349_io_x3; // @[MUL.scala 102:19]
  wire  m_2349_io_s; // @[MUL.scala 102:19]
  wire  m_2349_io_cout; // @[MUL.scala 102:19]
  wire  m_2350_io_x1; // @[MUL.scala 102:19]
  wire  m_2350_io_x2; // @[MUL.scala 102:19]
  wire  m_2350_io_x3; // @[MUL.scala 102:19]
  wire  m_2350_io_s; // @[MUL.scala 102:19]
  wire  m_2350_io_cout; // @[MUL.scala 102:19]
  wire  m_2351_io_x1; // @[MUL.scala 102:19]
  wire  m_2351_io_x2; // @[MUL.scala 102:19]
  wire  m_2351_io_x3; // @[MUL.scala 102:19]
  wire  m_2351_io_s; // @[MUL.scala 102:19]
  wire  m_2351_io_cout; // @[MUL.scala 102:19]
  wire  m_2352_io_x1; // @[MUL.scala 102:19]
  wire  m_2352_io_x2; // @[MUL.scala 102:19]
  wire  m_2352_io_x3; // @[MUL.scala 102:19]
  wire  m_2352_io_s; // @[MUL.scala 102:19]
  wire  m_2352_io_cout; // @[MUL.scala 102:19]
  wire  m_2353_io_x1; // @[MUL.scala 102:19]
  wire  m_2353_io_x2; // @[MUL.scala 102:19]
  wire  m_2353_io_x3; // @[MUL.scala 102:19]
  wire  m_2353_io_s; // @[MUL.scala 102:19]
  wire  m_2353_io_cout; // @[MUL.scala 102:19]
  wire  m_2354_io_x1; // @[MUL.scala 102:19]
  wire  m_2354_io_x2; // @[MUL.scala 102:19]
  wire  m_2354_io_x3; // @[MUL.scala 102:19]
  wire  m_2354_io_s; // @[MUL.scala 102:19]
  wire  m_2354_io_cout; // @[MUL.scala 102:19]
  wire  m_2355_io_x1; // @[MUL.scala 102:19]
  wire  m_2355_io_x2; // @[MUL.scala 102:19]
  wire  m_2355_io_x3; // @[MUL.scala 102:19]
  wire  m_2355_io_s; // @[MUL.scala 102:19]
  wire  m_2355_io_cout; // @[MUL.scala 102:19]
  wire  m_2356_io_x1; // @[MUL.scala 102:19]
  wire  m_2356_io_x2; // @[MUL.scala 102:19]
  wire  m_2356_io_x3; // @[MUL.scala 102:19]
  wire  m_2356_io_s; // @[MUL.scala 102:19]
  wire  m_2356_io_cout; // @[MUL.scala 102:19]
  wire  m_2357_io_x1; // @[MUL.scala 102:19]
  wire  m_2357_io_x2; // @[MUL.scala 102:19]
  wire  m_2357_io_x3; // @[MUL.scala 102:19]
  wire  m_2357_io_s; // @[MUL.scala 102:19]
  wire  m_2357_io_cout; // @[MUL.scala 102:19]
  wire  m_2358_io_x1; // @[MUL.scala 102:19]
  wire  m_2358_io_x2; // @[MUL.scala 102:19]
  wire  m_2358_io_x3; // @[MUL.scala 102:19]
  wire  m_2358_io_s; // @[MUL.scala 102:19]
  wire  m_2358_io_cout; // @[MUL.scala 102:19]
  wire  m_2359_io_x1; // @[MUL.scala 102:19]
  wire  m_2359_io_x2; // @[MUL.scala 102:19]
  wire  m_2359_io_x3; // @[MUL.scala 102:19]
  wire  m_2359_io_s; // @[MUL.scala 102:19]
  wire  m_2359_io_cout; // @[MUL.scala 102:19]
  wire  m_2360_io_x1; // @[MUL.scala 102:19]
  wire  m_2360_io_x2; // @[MUL.scala 102:19]
  wire  m_2360_io_x3; // @[MUL.scala 102:19]
  wire  m_2360_io_s; // @[MUL.scala 102:19]
  wire  m_2360_io_cout; // @[MUL.scala 102:19]
  wire  m_2361_io_x1; // @[MUL.scala 102:19]
  wire  m_2361_io_x2; // @[MUL.scala 102:19]
  wire  m_2361_io_x3; // @[MUL.scala 102:19]
  wire  m_2361_io_s; // @[MUL.scala 102:19]
  wire  m_2361_io_cout; // @[MUL.scala 102:19]
  wire  m_2362_io_x1; // @[MUL.scala 102:19]
  wire  m_2362_io_x2; // @[MUL.scala 102:19]
  wire  m_2362_io_x3; // @[MUL.scala 102:19]
  wire  m_2362_io_s; // @[MUL.scala 102:19]
  wire  m_2362_io_cout; // @[MUL.scala 102:19]
  wire  m_2363_io_x1; // @[MUL.scala 102:19]
  wire  m_2363_io_x2; // @[MUL.scala 102:19]
  wire  m_2363_io_x3; // @[MUL.scala 102:19]
  wire  m_2363_io_s; // @[MUL.scala 102:19]
  wire  m_2363_io_cout; // @[MUL.scala 102:19]
  wire  m_2364_io_x1; // @[MUL.scala 102:19]
  wire  m_2364_io_x2; // @[MUL.scala 102:19]
  wire  m_2364_io_x3; // @[MUL.scala 102:19]
  wire  m_2364_io_s; // @[MUL.scala 102:19]
  wire  m_2364_io_cout; // @[MUL.scala 102:19]
  wire  m_2365_io_x1; // @[MUL.scala 102:19]
  wire  m_2365_io_x2; // @[MUL.scala 102:19]
  wire  m_2365_io_x3; // @[MUL.scala 102:19]
  wire  m_2365_io_s; // @[MUL.scala 102:19]
  wire  m_2365_io_cout; // @[MUL.scala 102:19]
  wire  m_2366_io_x1; // @[MUL.scala 102:19]
  wire  m_2366_io_x2; // @[MUL.scala 102:19]
  wire  m_2366_io_x3; // @[MUL.scala 102:19]
  wire  m_2366_io_s; // @[MUL.scala 102:19]
  wire  m_2366_io_cout; // @[MUL.scala 102:19]
  wire  m_2367_io_x1; // @[MUL.scala 102:19]
  wire  m_2367_io_x2; // @[MUL.scala 102:19]
  wire  m_2367_io_x3; // @[MUL.scala 102:19]
  wire  m_2367_io_s; // @[MUL.scala 102:19]
  wire  m_2367_io_cout; // @[MUL.scala 102:19]
  wire  m_2368_io_x1; // @[MUL.scala 102:19]
  wire  m_2368_io_x2; // @[MUL.scala 102:19]
  wire  m_2368_io_x3; // @[MUL.scala 102:19]
  wire  m_2368_io_s; // @[MUL.scala 102:19]
  wire  m_2368_io_cout; // @[MUL.scala 102:19]
  wire  m_2369_io_x1; // @[MUL.scala 102:19]
  wire  m_2369_io_x2; // @[MUL.scala 102:19]
  wire  m_2369_io_x3; // @[MUL.scala 102:19]
  wire  m_2369_io_s; // @[MUL.scala 102:19]
  wire  m_2369_io_cout; // @[MUL.scala 102:19]
  wire  m_2370_io_x1; // @[MUL.scala 102:19]
  wire  m_2370_io_x2; // @[MUL.scala 102:19]
  wire  m_2370_io_x3; // @[MUL.scala 102:19]
  wire  m_2370_io_s; // @[MUL.scala 102:19]
  wire  m_2370_io_cout; // @[MUL.scala 102:19]
  wire  m_2371_io_x1; // @[MUL.scala 102:19]
  wire  m_2371_io_x2; // @[MUL.scala 102:19]
  wire  m_2371_io_x3; // @[MUL.scala 102:19]
  wire  m_2371_io_s; // @[MUL.scala 102:19]
  wire  m_2371_io_cout; // @[MUL.scala 102:19]
  wire  m_2372_io_x1; // @[MUL.scala 102:19]
  wire  m_2372_io_x2; // @[MUL.scala 102:19]
  wire  m_2372_io_x3; // @[MUL.scala 102:19]
  wire  m_2372_io_s; // @[MUL.scala 102:19]
  wire  m_2372_io_cout; // @[MUL.scala 102:19]
  wire  m_2373_io_x1; // @[MUL.scala 102:19]
  wire  m_2373_io_x2; // @[MUL.scala 102:19]
  wire  m_2373_io_x3; // @[MUL.scala 102:19]
  wire  m_2373_io_s; // @[MUL.scala 102:19]
  wire  m_2373_io_cout; // @[MUL.scala 102:19]
  wire  m_2374_io_x1; // @[MUL.scala 102:19]
  wire  m_2374_io_x2; // @[MUL.scala 102:19]
  wire  m_2374_io_x3; // @[MUL.scala 102:19]
  wire  m_2374_io_s; // @[MUL.scala 102:19]
  wire  m_2374_io_cout; // @[MUL.scala 102:19]
  wire  m_2375_io_x1; // @[MUL.scala 102:19]
  wire  m_2375_io_x2; // @[MUL.scala 102:19]
  wire  m_2375_io_x3; // @[MUL.scala 102:19]
  wire  m_2375_io_s; // @[MUL.scala 102:19]
  wire  m_2375_io_cout; // @[MUL.scala 102:19]
  wire  m_2376_io_x1; // @[MUL.scala 102:19]
  wire  m_2376_io_x2; // @[MUL.scala 102:19]
  wire  m_2376_io_x3; // @[MUL.scala 102:19]
  wire  m_2376_io_s; // @[MUL.scala 102:19]
  wire  m_2376_io_cout; // @[MUL.scala 102:19]
  wire  m_2377_io_in_0; // @[MUL.scala 124:19]
  wire  m_2377_io_in_1; // @[MUL.scala 124:19]
  wire  m_2377_io_out_0; // @[MUL.scala 124:19]
  wire  m_2377_io_out_1; // @[MUL.scala 124:19]
  wire  m_2378_io_in_0; // @[MUL.scala 124:19]
  wire  m_2378_io_in_1; // @[MUL.scala 124:19]
  wire  m_2378_io_out_0; // @[MUL.scala 124:19]
  wire  m_2378_io_out_1; // @[MUL.scala 124:19]
  wire  m_2379_io_in_0; // @[MUL.scala 124:19]
  wire  m_2379_io_in_1; // @[MUL.scala 124:19]
  wire  m_2379_io_out_0; // @[MUL.scala 124:19]
  wire  m_2379_io_out_1; // @[MUL.scala 124:19]
  wire  m_2380_io_in_0; // @[MUL.scala 124:19]
  wire  m_2380_io_in_1; // @[MUL.scala 124:19]
  wire  m_2380_io_out_0; // @[MUL.scala 124:19]
  wire  m_2380_io_out_1; // @[MUL.scala 124:19]
  wire  m_2381_io_in_0; // @[MUL.scala 124:19]
  wire  m_2381_io_in_1; // @[MUL.scala 124:19]
  wire  m_2381_io_out_0; // @[MUL.scala 124:19]
  wire  m_2381_io_out_1; // @[MUL.scala 124:19]
  wire  m_2382_io_in_0; // @[MUL.scala 124:19]
  wire  m_2382_io_in_1; // @[MUL.scala 124:19]
  wire  m_2382_io_out_0; // @[MUL.scala 124:19]
  wire  m_2382_io_out_1; // @[MUL.scala 124:19]
  wire  m_2383_io_in_0; // @[MUL.scala 124:19]
  wire  m_2383_io_in_1; // @[MUL.scala 124:19]
  wire  m_2383_io_out_0; // @[MUL.scala 124:19]
  wire  m_2383_io_out_1; // @[MUL.scala 124:19]
  wire  m_2384_io_in_0; // @[MUL.scala 124:19]
  wire  m_2384_io_in_1; // @[MUL.scala 124:19]
  wire  m_2384_io_out_0; // @[MUL.scala 124:19]
  wire  m_2384_io_out_1; // @[MUL.scala 124:19]
  wire  m_2385_io_in_0; // @[MUL.scala 124:19]
  wire  m_2385_io_in_1; // @[MUL.scala 124:19]
  wire  m_2385_io_out_0; // @[MUL.scala 124:19]
  wire  m_2385_io_out_1; // @[MUL.scala 124:19]
  wire  m_2386_io_in_0; // @[MUL.scala 124:19]
  wire  m_2386_io_in_1; // @[MUL.scala 124:19]
  wire  m_2386_io_out_0; // @[MUL.scala 124:19]
  wire  m_2386_io_out_1; // @[MUL.scala 124:19]
  wire  m_2387_io_in_0; // @[MUL.scala 124:19]
  wire  m_2387_io_in_1; // @[MUL.scala 124:19]
  wire  m_2387_io_out_0; // @[MUL.scala 124:19]
  wire  m_2387_io_out_1; // @[MUL.scala 124:19]
  wire  m_2388_io_in_0; // @[MUL.scala 124:19]
  wire  m_2388_io_in_1; // @[MUL.scala 124:19]
  wire  m_2388_io_out_0; // @[MUL.scala 124:19]
  wire  m_2388_io_out_1; // @[MUL.scala 124:19]
  wire  m_2389_io_in_0; // @[MUL.scala 124:19]
  wire  m_2389_io_in_1; // @[MUL.scala 124:19]
  wire  m_2389_io_out_0; // @[MUL.scala 124:19]
  wire  m_2389_io_out_1; // @[MUL.scala 124:19]
  wire  m_2390_io_in_0; // @[MUL.scala 124:19]
  wire  m_2390_io_in_1; // @[MUL.scala 124:19]
  wire  m_2390_io_out_0; // @[MUL.scala 124:19]
  wire  m_2390_io_out_1; // @[MUL.scala 124:19]
  wire  m_2391_io_in_0; // @[MUL.scala 124:19]
  wire  m_2391_io_in_1; // @[MUL.scala 124:19]
  wire  m_2391_io_out_0; // @[MUL.scala 124:19]
  wire  m_2391_io_out_1; // @[MUL.scala 124:19]
  wire  m_2392_io_in_0; // @[MUL.scala 124:19]
  wire  m_2392_io_in_1; // @[MUL.scala 124:19]
  wire  m_2392_io_out_0; // @[MUL.scala 124:19]
  wire  m_2392_io_out_1; // @[MUL.scala 124:19]
  wire  m_2393_io_in_0; // @[MUL.scala 124:19]
  wire  m_2393_io_in_1; // @[MUL.scala 124:19]
  wire  m_2393_io_out_0; // @[MUL.scala 124:19]
  wire  m_2393_io_out_1; // @[MUL.scala 124:19]
  wire  m_2394_io_in_0; // @[MUL.scala 124:19]
  wire  m_2394_io_in_1; // @[MUL.scala 124:19]
  wire  m_2394_io_out_0; // @[MUL.scala 124:19]
  wire  m_2394_io_out_1; // @[MUL.scala 124:19]
  wire  m_2395_io_in_0; // @[MUL.scala 124:19]
  wire  m_2395_io_in_1; // @[MUL.scala 124:19]
  wire  m_2395_io_out_0; // @[MUL.scala 124:19]
  wire  m_2395_io_out_1; // @[MUL.scala 124:19]
  wire  m_2396_io_in_0; // @[MUL.scala 124:19]
  wire  m_2396_io_in_1; // @[MUL.scala 124:19]
  wire  m_2396_io_out_0; // @[MUL.scala 124:19]
  wire  m_2396_io_out_1; // @[MUL.scala 124:19]
  wire  m_2397_io_in_0; // @[MUL.scala 124:19]
  wire  m_2397_io_in_1; // @[MUL.scala 124:19]
  wire  m_2397_io_out_0; // @[MUL.scala 124:19]
  wire  m_2397_io_out_1; // @[MUL.scala 124:19]
  wire  m_2398_io_in_0; // @[MUL.scala 124:19]
  wire  m_2398_io_in_1; // @[MUL.scala 124:19]
  wire  m_2398_io_out_0; // @[MUL.scala 124:19]
  wire  m_2398_io_out_1; // @[MUL.scala 124:19]
  wire  m_2399_io_in_0; // @[MUL.scala 124:19]
  wire  m_2399_io_in_1; // @[MUL.scala 124:19]
  wire  m_2399_io_out_0; // @[MUL.scala 124:19]
  wire  m_2399_io_out_1; // @[MUL.scala 124:19]
  wire  m_2400_io_in_0; // @[MUL.scala 124:19]
  wire  m_2400_io_in_1; // @[MUL.scala 124:19]
  wire  m_2400_io_out_0; // @[MUL.scala 124:19]
  wire  m_2400_io_out_1; // @[MUL.scala 124:19]
  wire  m_2401_io_in_0; // @[MUL.scala 124:19]
  wire  m_2401_io_in_1; // @[MUL.scala 124:19]
  wire  m_2401_io_out_0; // @[MUL.scala 124:19]
  wire  m_2401_io_out_1; // @[MUL.scala 124:19]
  wire  m_2402_io_in_0; // @[MUL.scala 124:19]
  wire  m_2402_io_in_1; // @[MUL.scala 124:19]
  wire  m_2402_io_out_0; // @[MUL.scala 124:19]
  wire  m_2402_io_out_1; // @[MUL.scala 124:19]
  wire  m_2403_io_in_0; // @[MUL.scala 124:19]
  wire  m_2403_io_in_1; // @[MUL.scala 124:19]
  wire  m_2403_io_out_0; // @[MUL.scala 124:19]
  wire  m_2403_io_out_1; // @[MUL.scala 124:19]
  wire  m_2404_io_in_0; // @[MUL.scala 124:19]
  wire  m_2404_io_in_1; // @[MUL.scala 124:19]
  wire  m_2404_io_out_0; // @[MUL.scala 124:19]
  wire  m_2404_io_out_1; // @[MUL.scala 124:19]
  wire  m_2405_io_in_0; // @[MUL.scala 124:19]
  wire  m_2405_io_in_1; // @[MUL.scala 124:19]
  wire  m_2405_io_out_0; // @[MUL.scala 124:19]
  wire  m_2405_io_out_1; // @[MUL.scala 124:19]
  wire  m_2406_io_in_0; // @[MUL.scala 124:19]
  wire  m_2406_io_in_1; // @[MUL.scala 124:19]
  wire  m_2406_io_out_0; // @[MUL.scala 124:19]
  wire  m_2406_io_out_1; // @[MUL.scala 124:19]
  wire  m_2407_io_in_0; // @[MUL.scala 124:19]
  wire  m_2407_io_in_1; // @[MUL.scala 124:19]
  wire  m_2407_io_out_0; // @[MUL.scala 124:19]
  wire  m_2407_io_out_1; // @[MUL.scala 124:19]
  wire  m_2408_io_in_0; // @[MUL.scala 124:19]
  wire  m_2408_io_in_1; // @[MUL.scala 124:19]
  wire  m_2408_io_out_0; // @[MUL.scala 124:19]
  wire  m_2408_io_out_1; // @[MUL.scala 124:19]
  wire  m_2409_io_in_0; // @[MUL.scala 124:19]
  wire  m_2409_io_in_1; // @[MUL.scala 124:19]
  wire  m_2409_io_out_0; // @[MUL.scala 124:19]
  wire  m_2409_io_out_1; // @[MUL.scala 124:19]
  wire  m_2410_io_in_0; // @[MUL.scala 124:19]
  wire  m_2410_io_in_1; // @[MUL.scala 124:19]
  wire  m_2410_io_out_0; // @[MUL.scala 124:19]
  wire  m_2410_io_out_1; // @[MUL.scala 124:19]
  wire  m_2411_io_in_0; // @[MUL.scala 124:19]
  wire  m_2411_io_in_1; // @[MUL.scala 124:19]
  wire  m_2411_io_out_0; // @[MUL.scala 124:19]
  wire  m_2411_io_out_1; // @[MUL.scala 124:19]
  wire  m_2412_io_in_0; // @[MUL.scala 124:19]
  wire  m_2412_io_in_1; // @[MUL.scala 124:19]
  wire  m_2412_io_out_0; // @[MUL.scala 124:19]
  wire  m_2412_io_out_1; // @[MUL.scala 124:19]
  wire  m_2413_io_in_0; // @[MUL.scala 124:19]
  wire  m_2413_io_in_1; // @[MUL.scala 124:19]
  wire  m_2413_io_out_0; // @[MUL.scala 124:19]
  wire  m_2413_io_out_1; // @[MUL.scala 124:19]
  wire  m_2414_io_in_0; // @[MUL.scala 124:19]
  wire  m_2414_io_in_1; // @[MUL.scala 124:19]
  wire  m_2414_io_out_0; // @[MUL.scala 124:19]
  wire  m_2414_io_out_1; // @[MUL.scala 124:19]
  wire  m_2415_io_in_0; // @[MUL.scala 124:19]
  wire  m_2415_io_in_1; // @[MUL.scala 124:19]
  wire  m_2415_io_out_0; // @[MUL.scala 124:19]
  wire  m_2415_io_out_1; // @[MUL.scala 124:19]
  wire  m_2416_io_in_0; // @[MUL.scala 124:19]
  wire  m_2416_io_in_1; // @[MUL.scala 124:19]
  wire  m_2416_io_out_0; // @[MUL.scala 124:19]
  wire  m_2416_io_out_1; // @[MUL.scala 124:19]
  wire  m_2417_io_in_0; // @[MUL.scala 124:19]
  wire  m_2417_io_in_1; // @[MUL.scala 124:19]
  wire  m_2417_io_out_0; // @[MUL.scala 124:19]
  wire  m_2417_io_out_1; // @[MUL.scala 124:19]
  wire  m_2418_io_in_0; // @[MUL.scala 124:19]
  wire  m_2418_io_in_1; // @[MUL.scala 124:19]
  wire  m_2418_io_out_0; // @[MUL.scala 124:19]
  wire  m_2418_io_out_1; // @[MUL.scala 124:19]
  wire  m_2419_io_in_0; // @[MUL.scala 124:19]
  wire  m_2419_io_in_1; // @[MUL.scala 124:19]
  wire  m_2419_io_out_0; // @[MUL.scala 124:19]
  wire  m_2419_io_out_1; // @[MUL.scala 124:19]
  wire  m_2420_io_in_0; // @[MUL.scala 124:19]
  wire  m_2420_io_in_1; // @[MUL.scala 124:19]
  wire  m_2420_io_out_0; // @[MUL.scala 124:19]
  wire  m_2420_io_out_1; // @[MUL.scala 124:19]
  wire  m_2421_io_in_0; // @[MUL.scala 124:19]
  wire  m_2421_io_in_1; // @[MUL.scala 124:19]
  wire  m_2421_io_out_0; // @[MUL.scala 124:19]
  wire  m_2421_io_out_1; // @[MUL.scala 124:19]
  wire  m_2422_io_in_0; // @[MUL.scala 124:19]
  wire  m_2422_io_in_1; // @[MUL.scala 124:19]
  wire  m_2422_io_out_0; // @[MUL.scala 124:19]
  wire  m_2422_io_out_1; // @[MUL.scala 124:19]
  wire  m_2423_io_in_0; // @[MUL.scala 124:19]
  wire  m_2423_io_in_1; // @[MUL.scala 124:19]
  wire  m_2423_io_out_0; // @[MUL.scala 124:19]
  wire  m_2423_io_out_1; // @[MUL.scala 124:19]
  wire  m_2424_io_in_0; // @[MUL.scala 124:19]
  wire  m_2424_io_in_1; // @[MUL.scala 124:19]
  wire  m_2424_io_out_0; // @[MUL.scala 124:19]
  wire  m_2424_io_out_1; // @[MUL.scala 124:19]
  wire  m_2425_io_in_0; // @[MUL.scala 124:19]
  wire  m_2425_io_in_1; // @[MUL.scala 124:19]
  wire  m_2425_io_out_0; // @[MUL.scala 124:19]
  wire  m_2425_io_out_1; // @[MUL.scala 124:19]
  wire  m_2426_io_in_0; // @[MUL.scala 124:19]
  wire  m_2426_io_in_1; // @[MUL.scala 124:19]
  wire  m_2426_io_out_0; // @[MUL.scala 124:19]
  wire  m_2426_io_out_1; // @[MUL.scala 124:19]
  wire  m_2427_io_in_0; // @[MUL.scala 124:19]
  wire  m_2427_io_in_1; // @[MUL.scala 124:19]
  wire  m_2427_io_out_0; // @[MUL.scala 124:19]
  wire  m_2427_io_out_1; // @[MUL.scala 124:19]
  wire  m_2428_io_in_0; // @[MUL.scala 124:19]
  wire  m_2428_io_in_1; // @[MUL.scala 124:19]
  wire  m_2428_io_out_0; // @[MUL.scala 124:19]
  wire  m_2428_io_out_1; // @[MUL.scala 124:19]
  wire  m_2429_io_in_0; // @[MUL.scala 124:19]
  wire  m_2429_io_in_1; // @[MUL.scala 124:19]
  wire  m_2429_io_out_0; // @[MUL.scala 124:19]
  wire  m_2429_io_out_1; // @[MUL.scala 124:19]
  wire  m_2430_io_in_0; // @[MUL.scala 124:19]
  wire  m_2430_io_in_1; // @[MUL.scala 124:19]
  wire  m_2430_io_out_0; // @[MUL.scala 124:19]
  wire  m_2430_io_out_1; // @[MUL.scala 124:19]
  wire  m_2431_io_in_0; // @[MUL.scala 124:19]
  wire  m_2431_io_in_1; // @[MUL.scala 124:19]
  wire  m_2431_io_out_0; // @[MUL.scala 124:19]
  wire  m_2431_io_out_1; // @[MUL.scala 124:19]
  wire  m_2432_io_in_0; // @[MUL.scala 124:19]
  wire  m_2432_io_in_1; // @[MUL.scala 124:19]
  wire  m_2432_io_out_0; // @[MUL.scala 124:19]
  wire  m_2432_io_out_1; // @[MUL.scala 124:19]
  wire  m_2433_io_in_0; // @[MUL.scala 124:19]
  wire  m_2433_io_in_1; // @[MUL.scala 124:19]
  wire  m_2433_io_out_0; // @[MUL.scala 124:19]
  wire  m_2433_io_out_1; // @[MUL.scala 124:19]
  wire  m_2434_io_in_0; // @[MUL.scala 124:19]
  wire  m_2434_io_in_1; // @[MUL.scala 124:19]
  wire  m_2434_io_out_0; // @[MUL.scala 124:19]
  wire  m_2434_io_out_1; // @[MUL.scala 124:19]
  wire  m_2435_io_in_0; // @[MUL.scala 124:19]
  wire  m_2435_io_in_1; // @[MUL.scala 124:19]
  wire  m_2435_io_out_0; // @[MUL.scala 124:19]
  wire  m_2435_io_out_1; // @[MUL.scala 124:19]
  wire  m_2436_io_in_0; // @[MUL.scala 124:19]
  wire  m_2436_io_in_1; // @[MUL.scala 124:19]
  wire  m_2436_io_out_0; // @[MUL.scala 124:19]
  wire  m_2436_io_out_1; // @[MUL.scala 124:19]
  wire  m_2437_io_in_0; // @[MUL.scala 124:19]
  wire  m_2437_io_in_1; // @[MUL.scala 124:19]
  wire  m_2437_io_out_0; // @[MUL.scala 124:19]
  wire  m_2437_io_out_1; // @[MUL.scala 124:19]
  wire  m_2438_io_in_0; // @[MUL.scala 124:19]
  wire  m_2438_io_in_1; // @[MUL.scala 124:19]
  wire  m_2438_io_out_0; // @[MUL.scala 124:19]
  wire  m_2438_io_out_1; // @[MUL.scala 124:19]
  wire  m_2439_io_in_0; // @[MUL.scala 124:19]
  wire  m_2439_io_in_1; // @[MUL.scala 124:19]
  wire  m_2439_io_out_0; // @[MUL.scala 124:19]
  wire  m_2439_io_out_1; // @[MUL.scala 124:19]
  wire  m_2440_io_in_0; // @[MUL.scala 124:19]
  wire  m_2440_io_in_1; // @[MUL.scala 124:19]
  wire  m_2440_io_out_0; // @[MUL.scala 124:19]
  wire  m_2440_io_out_1; // @[MUL.scala 124:19]
  wire  m_2441_io_in_0; // @[MUL.scala 124:19]
  wire  m_2441_io_in_1; // @[MUL.scala 124:19]
  wire  m_2441_io_out_0; // @[MUL.scala 124:19]
  wire  m_2441_io_out_1; // @[MUL.scala 124:19]
  wire  m_2442_io_in_0; // @[MUL.scala 124:19]
  wire  m_2442_io_in_1; // @[MUL.scala 124:19]
  wire  m_2442_io_out_0; // @[MUL.scala 124:19]
  wire  m_2442_io_out_1; // @[MUL.scala 124:19]
  wire  m_2443_io_in_0; // @[MUL.scala 124:19]
  wire  m_2443_io_in_1; // @[MUL.scala 124:19]
  wire  m_2443_io_out_0; // @[MUL.scala 124:19]
  wire  m_2443_io_out_1; // @[MUL.scala 124:19]
  wire  m_2444_io_in_0; // @[MUL.scala 124:19]
  wire  m_2444_io_in_1; // @[MUL.scala 124:19]
  wire  m_2444_io_out_0; // @[MUL.scala 124:19]
  wire  m_2444_io_out_1; // @[MUL.scala 124:19]
  wire  m_2445_io_in_0; // @[MUL.scala 124:19]
  wire  m_2445_io_in_1; // @[MUL.scala 124:19]
  wire  m_2445_io_out_0; // @[MUL.scala 124:19]
  wire  m_2445_io_out_1; // @[MUL.scala 124:19]
  wire  m_2446_io_in_0; // @[MUL.scala 124:19]
  wire  m_2446_io_in_1; // @[MUL.scala 124:19]
  wire  m_2446_io_out_0; // @[MUL.scala 124:19]
  wire  m_2446_io_out_1; // @[MUL.scala 124:19]
  wire  m_2447_io_in_0; // @[MUL.scala 124:19]
  wire  m_2447_io_in_1; // @[MUL.scala 124:19]
  wire  m_2447_io_out_0; // @[MUL.scala 124:19]
  wire  m_2447_io_out_1; // @[MUL.scala 124:19]
  wire  m_2448_io_in_0; // @[MUL.scala 124:19]
  wire  m_2448_io_in_1; // @[MUL.scala 124:19]
  wire  m_2448_io_out_0; // @[MUL.scala 124:19]
  wire  m_2448_io_out_1; // @[MUL.scala 124:19]
  wire  m_2449_io_in_0; // @[MUL.scala 124:19]
  wire  m_2449_io_in_1; // @[MUL.scala 124:19]
  wire  m_2449_io_out_0; // @[MUL.scala 124:19]
  wire  m_2449_io_out_1; // @[MUL.scala 124:19]
  wire  m_2450_io_in_0; // @[MUL.scala 124:19]
  wire  m_2450_io_in_1; // @[MUL.scala 124:19]
  wire  m_2450_io_out_0; // @[MUL.scala 124:19]
  wire  m_2450_io_out_1; // @[MUL.scala 124:19]
  wire  m_2451_io_in_0; // @[MUL.scala 124:19]
  wire  m_2451_io_in_1; // @[MUL.scala 124:19]
  wire  m_2451_io_out_0; // @[MUL.scala 124:19]
  wire  m_2451_io_out_1; // @[MUL.scala 124:19]
  wire  m_2452_io_in_0; // @[MUL.scala 124:19]
  wire  m_2452_io_in_1; // @[MUL.scala 124:19]
  wire  m_2452_io_out_0; // @[MUL.scala 124:19]
  wire  m_2452_io_out_1; // @[MUL.scala 124:19]
  wire  m_2453_io_in_0; // @[MUL.scala 124:19]
  wire  m_2453_io_in_1; // @[MUL.scala 124:19]
  wire  m_2453_io_out_0; // @[MUL.scala 124:19]
  wire  m_2453_io_out_1; // @[MUL.scala 124:19]
  wire  m_2454_io_in_0; // @[MUL.scala 124:19]
  wire  m_2454_io_in_1; // @[MUL.scala 124:19]
  wire  m_2454_io_out_0; // @[MUL.scala 124:19]
  wire  m_2454_io_out_1; // @[MUL.scala 124:19]
  wire  m_2455_io_in_0; // @[MUL.scala 124:19]
  wire  m_2455_io_in_1; // @[MUL.scala 124:19]
  wire  m_2455_io_out_0; // @[MUL.scala 124:19]
  wire  m_2455_io_out_1; // @[MUL.scala 124:19]
  wire  m_2456_io_in_0; // @[MUL.scala 124:19]
  wire  m_2456_io_in_1; // @[MUL.scala 124:19]
  wire  m_2456_io_out_0; // @[MUL.scala 124:19]
  wire  m_2456_io_out_1; // @[MUL.scala 124:19]
  wire  m_2457_io_in_0; // @[MUL.scala 124:19]
  wire  m_2457_io_in_1; // @[MUL.scala 124:19]
  wire  m_2457_io_out_0; // @[MUL.scala 124:19]
  wire  m_2457_io_out_1; // @[MUL.scala 124:19]
  wire  m_2458_io_in_0; // @[MUL.scala 124:19]
  wire  m_2458_io_in_1; // @[MUL.scala 124:19]
  wire  m_2458_io_out_0; // @[MUL.scala 124:19]
  wire  m_2458_io_out_1; // @[MUL.scala 124:19]
  wire  m_2459_io_in_0; // @[MUL.scala 124:19]
  wire  m_2459_io_in_1; // @[MUL.scala 124:19]
  wire  m_2459_io_out_0; // @[MUL.scala 124:19]
  wire  m_2459_io_out_1; // @[MUL.scala 124:19]
  wire  m_2460_io_in_0; // @[MUL.scala 124:19]
  wire  m_2460_io_in_1; // @[MUL.scala 124:19]
  wire  m_2460_io_out_0; // @[MUL.scala 124:19]
  wire  m_2460_io_out_1; // @[MUL.scala 124:19]
  wire  m_2461_io_in_0; // @[MUL.scala 124:19]
  wire  m_2461_io_in_1; // @[MUL.scala 124:19]
  wire  m_2461_io_out_0; // @[MUL.scala 124:19]
  wire  m_2461_io_out_1; // @[MUL.scala 124:19]
  wire  m_2462_io_x1; // @[MUL.scala 102:19]
  wire  m_2462_io_x2; // @[MUL.scala 102:19]
  wire  m_2462_io_x3; // @[MUL.scala 102:19]
  wire  m_2462_io_s; // @[MUL.scala 102:19]
  wire  m_2462_io_cout; // @[MUL.scala 102:19]
  wire  m_2463_io_x1; // @[MUL.scala 102:19]
  wire  m_2463_io_x2; // @[MUL.scala 102:19]
  wire  m_2463_io_x3; // @[MUL.scala 102:19]
  wire  m_2463_io_s; // @[MUL.scala 102:19]
  wire  m_2463_io_cout; // @[MUL.scala 102:19]
  wire  m_2464_io_x1; // @[MUL.scala 102:19]
  wire  m_2464_io_x2; // @[MUL.scala 102:19]
  wire  m_2464_io_x3; // @[MUL.scala 102:19]
  wire  m_2464_io_s; // @[MUL.scala 102:19]
  wire  m_2464_io_cout; // @[MUL.scala 102:19]
  wire  m_2465_io_x1; // @[MUL.scala 102:19]
  wire  m_2465_io_x2; // @[MUL.scala 102:19]
  wire  m_2465_io_x3; // @[MUL.scala 102:19]
  wire  m_2465_io_s; // @[MUL.scala 102:19]
  wire  m_2465_io_cout; // @[MUL.scala 102:19]
  wire  m_2466_io_x1; // @[MUL.scala 102:19]
  wire  m_2466_io_x2; // @[MUL.scala 102:19]
  wire  m_2466_io_x3; // @[MUL.scala 102:19]
  wire  m_2466_io_s; // @[MUL.scala 102:19]
  wire  m_2466_io_cout; // @[MUL.scala 102:19]
  wire  m_2467_io_x1; // @[MUL.scala 102:19]
  wire  m_2467_io_x2; // @[MUL.scala 102:19]
  wire  m_2467_io_x3; // @[MUL.scala 102:19]
  wire  m_2467_io_s; // @[MUL.scala 102:19]
  wire  m_2467_io_cout; // @[MUL.scala 102:19]
  wire  m_2468_io_x1; // @[MUL.scala 102:19]
  wire  m_2468_io_x2; // @[MUL.scala 102:19]
  wire  m_2468_io_x3; // @[MUL.scala 102:19]
  wire  m_2468_io_s; // @[MUL.scala 102:19]
  wire  m_2468_io_cout; // @[MUL.scala 102:19]
  wire  m_2469_io_x1; // @[MUL.scala 102:19]
  wire  m_2469_io_x2; // @[MUL.scala 102:19]
  wire  m_2469_io_x3; // @[MUL.scala 102:19]
  wire  m_2469_io_s; // @[MUL.scala 102:19]
  wire  m_2469_io_cout; // @[MUL.scala 102:19]
  wire  m_2470_io_x1; // @[MUL.scala 102:19]
  wire  m_2470_io_x2; // @[MUL.scala 102:19]
  wire  m_2470_io_x3; // @[MUL.scala 102:19]
  wire  m_2470_io_s; // @[MUL.scala 102:19]
  wire  m_2470_io_cout; // @[MUL.scala 102:19]
  wire  m_2471_io_x1; // @[MUL.scala 102:19]
  wire  m_2471_io_x2; // @[MUL.scala 102:19]
  wire  m_2471_io_x3; // @[MUL.scala 102:19]
  wire  m_2471_io_s; // @[MUL.scala 102:19]
  wire  m_2471_io_cout; // @[MUL.scala 102:19]
  wire  m_2472_io_x1; // @[MUL.scala 102:19]
  wire  m_2472_io_x2; // @[MUL.scala 102:19]
  wire  m_2472_io_x3; // @[MUL.scala 102:19]
  wire  m_2472_io_s; // @[MUL.scala 102:19]
  wire  m_2472_io_cout; // @[MUL.scala 102:19]
  wire  m_2473_io_x1; // @[MUL.scala 102:19]
  wire  m_2473_io_x2; // @[MUL.scala 102:19]
  wire  m_2473_io_x3; // @[MUL.scala 102:19]
  wire  m_2473_io_s; // @[MUL.scala 102:19]
  wire  m_2473_io_cout; // @[MUL.scala 102:19]
  wire  m_2474_io_x1; // @[MUL.scala 102:19]
  wire  m_2474_io_x2; // @[MUL.scala 102:19]
  wire  m_2474_io_x3; // @[MUL.scala 102:19]
  wire  m_2474_io_s; // @[MUL.scala 102:19]
  wire  m_2474_io_cout; // @[MUL.scala 102:19]
  wire  m_2475_io_x1; // @[MUL.scala 102:19]
  wire  m_2475_io_x2; // @[MUL.scala 102:19]
  wire  m_2475_io_x3; // @[MUL.scala 102:19]
  wire  m_2475_io_s; // @[MUL.scala 102:19]
  wire  m_2475_io_cout; // @[MUL.scala 102:19]
  wire  m_2476_io_x1; // @[MUL.scala 102:19]
  wire  m_2476_io_x2; // @[MUL.scala 102:19]
  wire  m_2476_io_x3; // @[MUL.scala 102:19]
  wire  m_2476_io_s; // @[MUL.scala 102:19]
  wire  m_2476_io_cout; // @[MUL.scala 102:19]
  wire  m_2477_io_x1; // @[MUL.scala 102:19]
  wire  m_2477_io_x2; // @[MUL.scala 102:19]
  wire  m_2477_io_x3; // @[MUL.scala 102:19]
  wire  m_2477_io_s; // @[MUL.scala 102:19]
  wire  m_2477_io_cout; // @[MUL.scala 102:19]
  wire  m_2478_io_x1; // @[MUL.scala 102:19]
  wire  m_2478_io_x2; // @[MUL.scala 102:19]
  wire  m_2478_io_x3; // @[MUL.scala 102:19]
  wire  m_2478_io_s; // @[MUL.scala 102:19]
  wire  m_2478_io_cout; // @[MUL.scala 102:19]
  wire  m_2479_io_x1; // @[MUL.scala 102:19]
  wire  m_2479_io_x2; // @[MUL.scala 102:19]
  wire  m_2479_io_x3; // @[MUL.scala 102:19]
  wire  m_2479_io_s; // @[MUL.scala 102:19]
  wire  m_2479_io_cout; // @[MUL.scala 102:19]
  wire  m_2480_io_x1; // @[MUL.scala 102:19]
  wire  m_2480_io_x2; // @[MUL.scala 102:19]
  wire  m_2480_io_x3; // @[MUL.scala 102:19]
  wire  m_2480_io_s; // @[MUL.scala 102:19]
  wire  m_2480_io_cout; // @[MUL.scala 102:19]
  wire  m_2481_io_x1; // @[MUL.scala 102:19]
  wire  m_2481_io_x2; // @[MUL.scala 102:19]
  wire  m_2481_io_x3; // @[MUL.scala 102:19]
  wire  m_2481_io_s; // @[MUL.scala 102:19]
  wire  m_2481_io_cout; // @[MUL.scala 102:19]
  wire  m_2482_io_x1; // @[MUL.scala 102:19]
  wire  m_2482_io_x2; // @[MUL.scala 102:19]
  wire  m_2482_io_x3; // @[MUL.scala 102:19]
  wire  m_2482_io_s; // @[MUL.scala 102:19]
  wire  m_2482_io_cout; // @[MUL.scala 102:19]
  wire  m_2483_io_in_0; // @[MUL.scala 124:19]
  wire  m_2483_io_in_1; // @[MUL.scala 124:19]
  wire  m_2483_io_out_0; // @[MUL.scala 124:19]
  wire  m_2483_io_out_1; // @[MUL.scala 124:19]
  wire  m_2484_io_in_0; // @[MUL.scala 124:19]
  wire  m_2484_io_in_1; // @[MUL.scala 124:19]
  wire  m_2484_io_out_0; // @[MUL.scala 124:19]
  wire  m_2484_io_out_1; // @[MUL.scala 124:19]
  wire  m_2485_io_in_0; // @[MUL.scala 124:19]
  wire  m_2485_io_in_1; // @[MUL.scala 124:19]
  wire  m_2485_io_out_0; // @[MUL.scala 124:19]
  wire  m_2485_io_out_1; // @[MUL.scala 124:19]
  wire  m_2486_io_in_0; // @[MUL.scala 124:19]
  wire  m_2486_io_in_1; // @[MUL.scala 124:19]
  wire  m_2486_io_out_0; // @[MUL.scala 124:19]
  wire  m_2486_io_out_1; // @[MUL.scala 124:19]
  wire  m_2487_io_in_0; // @[MUL.scala 124:19]
  wire  m_2487_io_in_1; // @[MUL.scala 124:19]
  wire  m_2487_io_out_0; // @[MUL.scala 124:19]
  wire  m_2487_io_out_1; // @[MUL.scala 124:19]
  wire  m_2488_io_in_0; // @[MUL.scala 124:19]
  wire  m_2488_io_in_1; // @[MUL.scala 124:19]
  wire  m_2488_io_out_0; // @[MUL.scala 124:19]
  wire  m_2488_io_out_1; // @[MUL.scala 124:19]
  wire  m_2489_io_in_0; // @[MUL.scala 124:19]
  wire  m_2489_io_in_1; // @[MUL.scala 124:19]
  wire  m_2489_io_out_0; // @[MUL.scala 124:19]
  wire  m_2489_io_out_1; // @[MUL.scala 124:19]
  wire  m_2490_io_in_0; // @[MUL.scala 124:19]
  wire  m_2490_io_in_1; // @[MUL.scala 124:19]
  wire  m_2490_io_out_0; // @[MUL.scala 124:19]
  wire  m_2490_io_out_1; // @[MUL.scala 124:19]
  wire  m_2491_io_in_0; // @[MUL.scala 124:19]
  wire  m_2491_io_in_1; // @[MUL.scala 124:19]
  wire  m_2491_io_out_0; // @[MUL.scala 124:19]
  wire  m_2491_io_out_1; // @[MUL.scala 124:19]
  wire  m_2492_io_in_0; // @[MUL.scala 124:19]
  wire  m_2492_io_in_1; // @[MUL.scala 124:19]
  wire  m_2492_io_out_0; // @[MUL.scala 124:19]
  wire  m_2492_io_out_1; // @[MUL.scala 124:19]
  wire  m_2493_io_in_0; // @[MUL.scala 124:19]
  wire  m_2493_io_in_1; // @[MUL.scala 124:19]
  wire  m_2493_io_out_0; // @[MUL.scala 124:19]
  wire  m_2493_io_out_1; // @[MUL.scala 124:19]
  wire  m_2494_io_in_0; // @[MUL.scala 124:19]
  wire  m_2494_io_in_1; // @[MUL.scala 124:19]
  wire  m_2494_io_out_0; // @[MUL.scala 124:19]
  wire  m_2494_io_out_1; // @[MUL.scala 124:19]
  wire  m_2495_io_in_0; // @[MUL.scala 124:19]
  wire  m_2495_io_in_1; // @[MUL.scala 124:19]
  wire  m_2495_io_out_0; // @[MUL.scala 124:19]
  wire  m_2495_io_out_1; // @[MUL.scala 124:19]
  wire  m_2496_io_in_0; // @[MUL.scala 124:19]
  wire  m_2496_io_in_1; // @[MUL.scala 124:19]
  wire  m_2496_io_out_0; // @[MUL.scala 124:19]
  wire  m_2496_io_out_1; // @[MUL.scala 124:19]
  wire  m_2497_io_in_0; // @[MUL.scala 124:19]
  wire  m_2497_io_in_1; // @[MUL.scala 124:19]
  wire  m_2497_io_out_0; // @[MUL.scala 124:19]
  wire  m_2497_io_out_1; // @[MUL.scala 124:19]
  wire  m_2498_io_in_0; // @[MUL.scala 124:19]
  wire  m_2498_io_in_1; // @[MUL.scala 124:19]
  wire  m_2498_io_out_0; // @[MUL.scala 124:19]
  wire  m_2498_io_out_1; // @[MUL.scala 124:19]
  wire  m_2499_io_in_0; // @[MUL.scala 124:19]
  wire  m_2499_io_in_1; // @[MUL.scala 124:19]
  wire  m_2499_io_out_0; // @[MUL.scala 124:19]
  wire  m_2499_io_out_1; // @[MUL.scala 124:19]
  wire  m_2500_io_in_0; // @[MUL.scala 124:19]
  wire  m_2500_io_in_1; // @[MUL.scala 124:19]
  wire  m_2500_io_out_0; // @[MUL.scala 124:19]
  wire  m_2500_io_out_1; // @[MUL.scala 124:19]
  wire  m_2501_io_in_0; // @[MUL.scala 124:19]
  wire  m_2501_io_in_1; // @[MUL.scala 124:19]
  wire  m_2501_io_out_0; // @[MUL.scala 124:19]
  wire  m_2501_io_out_1; // @[MUL.scala 124:19]
  wire  m_2502_io_in_0; // @[MUL.scala 124:19]
  wire  m_2502_io_in_1; // @[MUL.scala 124:19]
  wire  m_2502_io_out_0; // @[MUL.scala 124:19]
  wire  m_2502_io_out_1; // @[MUL.scala 124:19]
  wire  m_2503_io_in_0; // @[MUL.scala 124:19]
  wire  m_2503_io_in_1; // @[MUL.scala 124:19]
  wire  m_2503_io_out_0; // @[MUL.scala 124:19]
  wire  m_2503_io_out_1; // @[MUL.scala 124:19]
  wire  m_2504_io_in_0; // @[MUL.scala 124:19]
  wire  m_2504_io_in_1; // @[MUL.scala 124:19]
  wire  m_2504_io_out_0; // @[MUL.scala 124:19]
  wire  m_2504_io_out_1; // @[MUL.scala 124:19]
  wire  m_2505_io_in_0; // @[MUL.scala 124:19]
  wire  m_2505_io_in_1; // @[MUL.scala 124:19]
  wire  m_2505_io_out_0; // @[MUL.scala 124:19]
  wire  m_2505_io_out_1; // @[MUL.scala 124:19]
  wire  m_2506_io_in_0; // @[MUL.scala 124:19]
  wire  m_2506_io_in_1; // @[MUL.scala 124:19]
  wire  m_2506_io_out_0; // @[MUL.scala 124:19]
  wire  m_2506_io_out_1; // @[MUL.scala 124:19]
  wire  m_2507_io_in_0; // @[MUL.scala 124:19]
  wire  m_2507_io_in_1; // @[MUL.scala 124:19]
  wire  m_2507_io_out_0; // @[MUL.scala 124:19]
  wire  m_2507_io_out_1; // @[MUL.scala 124:19]
  wire  m_2508_io_in_0; // @[MUL.scala 124:19]
  wire  m_2508_io_in_1; // @[MUL.scala 124:19]
  wire  m_2508_io_out_0; // @[MUL.scala 124:19]
  wire  m_2508_io_out_1; // @[MUL.scala 124:19]
  wire  m_2509_io_in_0; // @[MUL.scala 124:19]
  wire  m_2509_io_in_1; // @[MUL.scala 124:19]
  wire  m_2509_io_out_0; // @[MUL.scala 124:19]
  wire  m_2509_io_out_1; // @[MUL.scala 124:19]
  wire  m_2510_io_in_0; // @[MUL.scala 124:19]
  wire  m_2510_io_in_1; // @[MUL.scala 124:19]
  wire  m_2510_io_out_0; // @[MUL.scala 124:19]
  wire  m_2510_io_out_1; // @[MUL.scala 124:19]
  wire  m_2511_io_in_0; // @[MUL.scala 124:19]
  wire  m_2511_io_in_1; // @[MUL.scala 124:19]
  wire  m_2511_io_out_0; // @[MUL.scala 124:19]
  wire  m_2511_io_out_1; // @[MUL.scala 124:19]
  wire  m_2512_io_in_0; // @[MUL.scala 124:19]
  wire  m_2512_io_in_1; // @[MUL.scala 124:19]
  wire  m_2512_io_out_0; // @[MUL.scala 124:19]
  wire  m_2512_io_out_1; // @[MUL.scala 124:19]
  wire  m_2513_io_in_0; // @[MUL.scala 124:19]
  wire  m_2513_io_in_1; // @[MUL.scala 124:19]
  wire  m_2513_io_out_0; // @[MUL.scala 124:19]
  wire  m_2513_io_out_1; // @[MUL.scala 124:19]
  wire  m_2514_io_in_0; // @[MUL.scala 124:19]
  wire  m_2514_io_in_1; // @[MUL.scala 124:19]
  wire  m_2514_io_out_0; // @[MUL.scala 124:19]
  wire  m_2514_io_out_1; // @[MUL.scala 124:19]
  wire  m_2515_io_in_0; // @[MUL.scala 124:19]
  wire  m_2515_io_in_1; // @[MUL.scala 124:19]
  wire  m_2515_io_out_0; // @[MUL.scala 124:19]
  wire  m_2515_io_out_1; // @[MUL.scala 124:19]
  wire  m_2516_io_in_0; // @[MUL.scala 124:19]
  wire  m_2516_io_in_1; // @[MUL.scala 124:19]
  wire  m_2516_io_out_0; // @[MUL.scala 124:19]
  wire  m_2516_io_out_1; // @[MUL.scala 124:19]
  wire  m_2517_io_in_0; // @[MUL.scala 124:19]
  wire  m_2517_io_in_1; // @[MUL.scala 124:19]
  wire  m_2517_io_out_0; // @[MUL.scala 124:19]
  wire  m_2517_io_out_1; // @[MUL.scala 124:19]
  wire  m_2518_io_in_0; // @[MUL.scala 124:19]
  wire  m_2518_io_in_1; // @[MUL.scala 124:19]
  wire  m_2518_io_out_0; // @[MUL.scala 124:19]
  wire  m_2518_io_out_1; // @[MUL.scala 124:19]
  wire  m_2519_io_in_0; // @[MUL.scala 124:19]
  wire  m_2519_io_in_1; // @[MUL.scala 124:19]
  wire  m_2519_io_out_0; // @[MUL.scala 124:19]
  wire  m_2519_io_out_1; // @[MUL.scala 124:19]
  wire  m_2520_io_in_0; // @[MUL.scala 124:19]
  wire  m_2520_io_in_1; // @[MUL.scala 124:19]
  wire  m_2520_io_out_0; // @[MUL.scala 124:19]
  wire  m_2520_io_out_1; // @[MUL.scala 124:19]
  wire  m_2521_io_in_0; // @[MUL.scala 124:19]
  wire  m_2521_io_in_1; // @[MUL.scala 124:19]
  wire  m_2521_io_out_0; // @[MUL.scala 124:19]
  wire  m_2521_io_out_1; // @[MUL.scala 124:19]
  wire  m_2522_io_in_0; // @[MUL.scala 124:19]
  wire  m_2522_io_in_1; // @[MUL.scala 124:19]
  wire  m_2522_io_out_0; // @[MUL.scala 124:19]
  wire  m_2522_io_out_1; // @[MUL.scala 124:19]
  wire  m_2523_io_in_0; // @[MUL.scala 124:19]
  wire  m_2523_io_in_1; // @[MUL.scala 124:19]
  wire  m_2523_io_out_0; // @[MUL.scala 124:19]
  wire  m_2523_io_out_1; // @[MUL.scala 124:19]
  wire  m_2524_io_in_0; // @[MUL.scala 124:19]
  wire  m_2524_io_in_1; // @[MUL.scala 124:19]
  wire  m_2524_io_out_0; // @[MUL.scala 124:19]
  wire  m_2524_io_out_1; // @[MUL.scala 124:19]
  wire  m_2525_io_in_0; // @[MUL.scala 124:19]
  wire  m_2525_io_in_1; // @[MUL.scala 124:19]
  wire  m_2525_io_out_0; // @[MUL.scala 124:19]
  wire  m_2525_io_out_1; // @[MUL.scala 124:19]
  wire  m_2526_io_in_0; // @[MUL.scala 124:19]
  wire  m_2526_io_in_1; // @[MUL.scala 124:19]
  wire  m_2526_io_out_0; // @[MUL.scala 124:19]
  wire  m_2526_io_out_1; // @[MUL.scala 124:19]
  wire  m_2527_io_in_0; // @[MUL.scala 124:19]
  wire  m_2527_io_in_1; // @[MUL.scala 124:19]
  wire  m_2527_io_out_0; // @[MUL.scala 124:19]
  wire  m_2527_io_out_1; // @[MUL.scala 124:19]
  wire  m_2528_io_in_0; // @[MUL.scala 124:19]
  wire  m_2528_io_in_1; // @[MUL.scala 124:19]
  wire  m_2528_io_out_0; // @[MUL.scala 124:19]
  wire  m_2528_io_out_1; // @[MUL.scala 124:19]
  wire  m_2529_io_in_0; // @[MUL.scala 124:19]
  wire  m_2529_io_in_1; // @[MUL.scala 124:19]
  wire  m_2529_io_out_0; // @[MUL.scala 124:19]
  wire  m_2529_io_out_1; // @[MUL.scala 124:19]
  wire  m_2530_io_in_0; // @[MUL.scala 124:19]
  wire  m_2530_io_in_1; // @[MUL.scala 124:19]
  wire  m_2530_io_out_0; // @[MUL.scala 124:19]
  wire  m_2530_io_out_1; // @[MUL.scala 124:19]
  wire  m_2531_io_in_0; // @[MUL.scala 124:19]
  wire  m_2531_io_in_1; // @[MUL.scala 124:19]
  wire  m_2531_io_out_0; // @[MUL.scala 124:19]
  wire  m_2531_io_out_1; // @[MUL.scala 124:19]
  wire  m_2532_io_in_0; // @[MUL.scala 124:19]
  wire  m_2532_io_in_1; // @[MUL.scala 124:19]
  wire  m_2532_io_out_0; // @[MUL.scala 124:19]
  wire  m_2532_io_out_1; // @[MUL.scala 124:19]
  wire  m_2533_io_in_0; // @[MUL.scala 124:19]
  wire  m_2533_io_in_1; // @[MUL.scala 124:19]
  wire  m_2533_io_out_0; // @[MUL.scala 124:19]
  wire  m_2533_io_out_1; // @[MUL.scala 124:19]
  wire  m_2534_io_in_0; // @[MUL.scala 124:19]
  wire  m_2534_io_in_1; // @[MUL.scala 124:19]
  wire  m_2534_io_out_0; // @[MUL.scala 124:19]
  wire  m_2534_io_out_1; // @[MUL.scala 124:19]
  wire [66:0] src1 = {2'h0,io_in_bits_ctrl_data_src1,1'h0}; // @[Cat.scala 31:58]
  wire  _T_88 = ~m_io_p[65]; // @[MUL.scala 313:93]
  wire  _T_157 = ~m_1_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_228 = ~m_2_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_299 = ~m_3_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_370 = ~m_4_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_441 = ~m_5_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_512 = ~m_6_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_583 = ~m_7_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_654 = ~m_8_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_725 = ~m_9_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_796 = ~m_10_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_867 = ~m_11_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_938 = ~m_12_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_1009 = ~m_13_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_1080 = ~m_14_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_1151 = ~m_15_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_1222 = ~m_16_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_1293 = ~m_17_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_1364 = ~m_18_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_1435 = ~m_19_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_1506 = ~m_20_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_1577 = ~m_21_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_1648 = ~m_22_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_1719 = ~m_23_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_1790 = ~m_24_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_1861 = ~m_25_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_1932 = ~m_26_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_2003 = ~m_27_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_2074 = ~m_28_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_2145 = ~m_29_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_2216 = ~m_30_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_2287 = ~m_31_io_p[65]; // @[MUL.scala 307:92]
  wire  _T_2358 = ~m_32_io_p[65]; // @[MUL.scala 316:92]
  reg  r; // @[Reg.scala 16:16]
  reg  r_1; // @[Reg.scala 16:16]
  reg  r_2; // @[Reg.scala 16:16]
  reg  r_3; // @[Reg.scala 16:16]
  reg  r_4; // @[Reg.scala 16:16]
  reg  r_5; // @[Reg.scala 16:16]
  reg  r_6; // @[Reg.scala 16:16]
  reg  r_7; // @[Reg.scala 16:16]
  reg  r_8; // @[Reg.scala 16:16]
  reg  r_9; // @[Reg.scala 16:16]
  reg  r_10; // @[Reg.scala 16:16]
  reg  r_11; // @[Reg.scala 16:16]
  reg  r_12; // @[Reg.scala 16:16]
  reg  r_13; // @[Reg.scala 16:16]
  reg  r_14; // @[Reg.scala 16:16]
  reg  r_15; // @[Reg.scala 16:16]
  reg  r_16; // @[Reg.scala 16:16]
  reg  r_17; // @[Reg.scala 16:16]
  reg  r_18; // @[Reg.scala 16:16]
  reg  r_19; // @[Reg.scala 16:16]
  reg  r_20; // @[Reg.scala 16:16]
  reg  r_21; // @[Reg.scala 16:16]
  reg  r_22; // @[Reg.scala 16:16]
  reg  r_23; // @[Reg.scala 16:16]
  reg  r_24; // @[Reg.scala 16:16]
  reg  r_25; // @[Reg.scala 16:16]
  reg  r_26; // @[Reg.scala 16:16]
  reg  r_27; // @[Reg.scala 16:16]
  reg  r_28; // @[Reg.scala 16:16]
  reg  r_29; // @[Reg.scala 16:16]
  reg  r_30; // @[Reg.scala 16:16]
  reg  r_31; // @[Reg.scala 16:16]
  reg  r_32; // @[Reg.scala 16:16]
  reg  r_33; // @[Reg.scala 16:16]
  reg  r_34; // @[Reg.scala 16:16]
  reg  r_35; // @[Reg.scala 16:16]
  reg  r_36; // @[Reg.scala 16:16]
  reg  r_37; // @[Reg.scala 16:16]
  reg  r_38; // @[Reg.scala 16:16]
  reg  r_39; // @[Reg.scala 16:16]
  reg  r_40; // @[Reg.scala 16:16]
  reg  r_41; // @[Reg.scala 16:16]
  reg  r_42; // @[Reg.scala 16:16]
  reg  r_43; // @[Reg.scala 16:16]
  reg  r_44; // @[Reg.scala 16:16]
  reg  r_45; // @[Reg.scala 16:16]
  reg  r_46; // @[Reg.scala 16:16]
  reg  r_47; // @[Reg.scala 16:16]
  reg  r_48; // @[Reg.scala 16:16]
  reg  r_49; // @[Reg.scala 16:16]
  reg  r_50; // @[Reg.scala 16:16]
  reg  r_51; // @[Reg.scala 16:16]
  reg  r_52; // @[Reg.scala 16:16]
  reg  r_53; // @[Reg.scala 16:16]
  reg  r_54; // @[Reg.scala 16:16]
  reg  r_55; // @[Reg.scala 16:16]
  reg  r_56; // @[Reg.scala 16:16]
  reg  r_57; // @[Reg.scala 16:16]
  reg  r_58; // @[Reg.scala 16:16]
  reg  r_59; // @[Reg.scala 16:16]
  reg  r_60; // @[Reg.scala 16:16]
  reg  r_61; // @[Reg.scala 16:16]
  reg  r_62; // @[Reg.scala 16:16]
  reg  r_63; // @[Reg.scala 16:16]
  reg  r_64; // @[Reg.scala 16:16]
  reg  r_65; // @[Reg.scala 16:16]
  reg  r_66; // @[Reg.scala 16:16]
  reg  r_67; // @[Reg.scala 16:16]
  reg  r_68; // @[Reg.scala 16:16]
  reg  r_69; // @[Reg.scala 16:16]
  reg  r_70; // @[Reg.scala 16:16]
  reg  r_71; // @[Reg.scala 16:16]
  reg  r_72; // @[Reg.scala 16:16]
  reg  r_73; // @[Reg.scala 16:16]
  reg  r_74; // @[Reg.scala 16:16]
  reg  r_75; // @[Reg.scala 16:16]
  reg  r_76; // @[Reg.scala 16:16]
  reg  r_77; // @[Reg.scala 16:16]
  reg  r_78; // @[Reg.scala 16:16]
  reg  r_79; // @[Reg.scala 16:16]
  reg  r_80; // @[Reg.scala 16:16]
  reg  r_81; // @[Reg.scala 16:16]
  reg  r_82; // @[Reg.scala 16:16]
  reg  r_83; // @[Reg.scala 16:16]
  reg  r_84; // @[Reg.scala 16:16]
  reg  r_85; // @[Reg.scala 16:16]
  reg  r_86; // @[Reg.scala 16:16]
  reg  r_87; // @[Reg.scala 16:16]
  reg  r_88; // @[Reg.scala 16:16]
  reg  r_89; // @[Reg.scala 16:16]
  reg  r_90; // @[Reg.scala 16:16]
  reg  r_91; // @[Reg.scala 16:16]
  reg  r_92; // @[Reg.scala 16:16]
  reg  r_93; // @[Reg.scala 16:16]
  reg  r_94; // @[Reg.scala 16:16]
  reg  r_95; // @[Reg.scala 16:16]
  reg  r_96; // @[Reg.scala 16:16]
  reg  r_97; // @[Reg.scala 16:16]
  reg  r_98; // @[Reg.scala 16:16]
  reg  r_99; // @[Reg.scala 16:16]
  reg  r_100; // @[Reg.scala 16:16]
  reg  r_101; // @[Reg.scala 16:16]
  reg  r_102; // @[Reg.scala 16:16]
  reg  r_103; // @[Reg.scala 16:16]
  reg  r_104; // @[Reg.scala 16:16]
  reg  r_105; // @[Reg.scala 16:16]
  reg  r_106; // @[Reg.scala 16:16]
  reg  r_107; // @[Reg.scala 16:16]
  reg  r_108; // @[Reg.scala 16:16]
  reg  r_109; // @[Reg.scala 16:16]
  reg  r_110; // @[Reg.scala 16:16]
  reg  r_111; // @[Reg.scala 16:16]
  reg  r_112; // @[Reg.scala 16:16]
  reg  r_113; // @[Reg.scala 16:16]
  reg  r_114; // @[Reg.scala 16:16]
  reg  r_115; // @[Reg.scala 16:16]
  reg  r_116; // @[Reg.scala 16:16]
  reg  r_117; // @[Reg.scala 16:16]
  reg  r_118; // @[Reg.scala 16:16]
  reg  r_119; // @[Reg.scala 16:16]
  reg  r_120; // @[Reg.scala 16:16]
  reg  r_121; // @[Reg.scala 16:16]
  reg  r_122; // @[Reg.scala 16:16]
  reg  r_123; // @[Reg.scala 16:16]
  reg  r_124; // @[Reg.scala 16:16]
  reg  r_125; // @[Reg.scala 16:16]
  reg  r_126; // @[Reg.scala 16:16]
  reg  r_127; // @[Reg.scala 16:16]
  reg  r_128; // @[Reg.scala 16:16]
  reg  r_129; // @[Reg.scala 16:16]
  reg  r_130; // @[Reg.scala 16:16]
  reg  r_131; // @[Reg.scala 16:16]
  reg  r_132; // @[Reg.scala 16:16]
  reg  r_133; // @[Reg.scala 16:16]
  reg  r_134; // @[Reg.scala 16:16]
  reg  r_135; // @[Reg.scala 16:16]
  reg  r_136; // @[Reg.scala 16:16]
  reg  r_137; // @[Reg.scala 16:16]
  reg  r_138; // @[Reg.scala 16:16]
  reg  r_139; // @[Reg.scala 16:16]
  reg  r_140; // @[Reg.scala 16:16]
  reg  r_141; // @[Reg.scala 16:16]
  reg  r_142; // @[Reg.scala 16:16]
  reg  r_143; // @[Reg.scala 16:16]
  reg  r_144; // @[Reg.scala 16:16]
  reg  r_145; // @[Reg.scala 16:16]
  reg  r_146; // @[Reg.scala 16:16]
  reg  r_147; // @[Reg.scala 16:16]
  reg  r_148; // @[Reg.scala 16:16]
  reg  r_149; // @[Reg.scala 16:16]
  reg  r_150; // @[Reg.scala 16:16]
  reg  r_151; // @[Reg.scala 16:16]
  reg  r_152; // @[Reg.scala 16:16]
  reg  r_153; // @[Reg.scala 16:16]
  reg  r_154; // @[Reg.scala 16:16]
  reg  r_155; // @[Reg.scala 16:16]
  reg  r_156; // @[Reg.scala 16:16]
  reg  r_157; // @[Reg.scala 16:16]
  reg  r_158; // @[Reg.scala 16:16]
  reg  r_159; // @[Reg.scala 16:16]
  reg  r_160; // @[Reg.scala 16:16]
  reg  r_161; // @[Reg.scala 16:16]
  reg  r_162; // @[Reg.scala 16:16]
  reg  r_163; // @[Reg.scala 16:16]
  reg  r_164; // @[Reg.scala 16:16]
  reg  r_165; // @[Reg.scala 16:16]
  reg  r_166; // @[Reg.scala 16:16]
  reg  r_167; // @[Reg.scala 16:16]
  reg  r_168; // @[Reg.scala 16:16]
  reg  r_169; // @[Reg.scala 16:16]
  reg  r_170; // @[Reg.scala 16:16]
  reg  r_171; // @[Reg.scala 16:16]
  reg  r_172; // @[Reg.scala 16:16]
  reg  r_173; // @[Reg.scala 16:16]
  reg  r_174; // @[Reg.scala 16:16]
  reg  r_175; // @[Reg.scala 16:16]
  reg  r_176; // @[Reg.scala 16:16]
  reg  r_177; // @[Reg.scala 16:16]
  reg  r_178; // @[Reg.scala 16:16]
  reg  r_179; // @[Reg.scala 16:16]
  reg  r_180; // @[Reg.scala 16:16]
  reg  r_181; // @[Reg.scala 16:16]
  reg  r_182; // @[Reg.scala 16:16]
  reg  r_183; // @[Reg.scala 16:16]
  reg  r_184; // @[Reg.scala 16:16]
  reg  r_185; // @[Reg.scala 16:16]
  reg  r_186; // @[Reg.scala 16:16]
  reg  r_187; // @[Reg.scala 16:16]
  reg  r_188; // @[Reg.scala 16:16]
  reg  r_189; // @[Reg.scala 16:16]
  reg  r_190; // @[Reg.scala 16:16]
  reg  r_191; // @[Reg.scala 16:16]
  reg  r_192; // @[Reg.scala 16:16]
  reg  r_193; // @[Reg.scala 16:16]
  reg  r_194; // @[Reg.scala 16:16]
  reg  r_195; // @[Reg.scala 16:16]
  reg  r_196; // @[Reg.scala 16:16]
  reg  r_197; // @[Reg.scala 16:16]
  reg  r_198; // @[Reg.scala 16:16]
  reg  r_199; // @[Reg.scala 16:16]
  reg  r_200; // @[Reg.scala 16:16]
  reg  r_201; // @[Reg.scala 16:16]
  reg  r_202; // @[Reg.scala 16:16]
  reg  r_203; // @[Reg.scala 16:16]
  reg  r_204; // @[Reg.scala 16:16]
  reg  r_205; // @[Reg.scala 16:16]
  reg  r_206; // @[Reg.scala 16:16]
  reg  r_207; // @[Reg.scala 16:16]
  reg  r_208; // @[Reg.scala 16:16]
  reg  r_209; // @[Reg.scala 16:16]
  reg  r_210; // @[Reg.scala 16:16]
  reg  r_211; // @[Reg.scala 16:16]
  reg  r_212; // @[Reg.scala 16:16]
  reg  r_213; // @[Reg.scala 16:16]
  reg  r_214; // @[Reg.scala 16:16]
  reg  r_215; // @[Reg.scala 16:16]
  reg  r_216; // @[Reg.scala 16:16]
  reg  r_217; // @[Reg.scala 16:16]
  reg  r_218; // @[Reg.scala 16:16]
  reg  r_219; // @[Reg.scala 16:16]
  reg  r_220; // @[Reg.scala 16:16]
  reg  r_221; // @[Reg.scala 16:16]
  reg  r_222; // @[Reg.scala 16:16]
  reg  r_223; // @[Reg.scala 16:16]
  reg  r_224; // @[Reg.scala 16:16]
  reg  r_225; // @[Reg.scala 16:16]
  reg  r_226; // @[Reg.scala 16:16]
  reg  r_227; // @[Reg.scala 16:16]
  reg  r_228; // @[Reg.scala 16:16]
  reg  r_229; // @[Reg.scala 16:16]
  reg  r_230; // @[Reg.scala 16:16]
  reg  r_231; // @[Reg.scala 16:16]
  reg  r_232; // @[Reg.scala 16:16]
  reg  r_233; // @[Reg.scala 16:16]
  reg  r_234; // @[Reg.scala 16:16]
  reg  r_235; // @[Reg.scala 16:16]
  reg  r_236; // @[Reg.scala 16:16]
  reg  r_237; // @[Reg.scala 16:16]
  reg  r_238; // @[Reg.scala 16:16]
  reg  r_239; // @[Reg.scala 16:16]
  reg  r_240; // @[Reg.scala 16:16]
  reg  r_241; // @[Reg.scala 16:16]
  reg  r_242; // @[Reg.scala 16:16]
  reg  r_243; // @[Reg.scala 16:16]
  reg  r_244; // @[Reg.scala 16:16]
  reg  r_245; // @[Reg.scala 16:16]
  reg  r_246; // @[Reg.scala 16:16]
  reg  r_247; // @[Reg.scala 16:16]
  reg  r_248; // @[Reg.scala 16:16]
  reg  r_249; // @[Reg.scala 16:16]
  reg  r_250; // @[Reg.scala 16:16]
  reg  r_251; // @[Reg.scala 16:16]
  reg  r_252; // @[Reg.scala 16:16]
  reg  r_253; // @[Reg.scala 16:16]
  reg  r_254; // @[Reg.scala 16:16]
  reg  r_255; // @[Reg.scala 16:16]
  reg  r_256; // @[Reg.scala 16:16]
  reg  r_257; // @[Reg.scala 16:16]
  reg  r_258; // @[Reg.scala 16:16]
  reg  r_259; // @[Reg.scala 16:16]
  reg  r_260; // @[Reg.scala 16:16]
  reg  r_261; // @[Reg.scala 16:16]
  reg  r_262; // @[Reg.scala 16:16]
  reg  r_263; // @[Reg.scala 16:16]
  reg  r_264; // @[Reg.scala 16:16]
  reg  r_265; // @[Reg.scala 16:16]
  reg  r_266; // @[Reg.scala 16:16]
  reg  r_267; // @[Reg.scala 16:16]
  reg  r_268; // @[Reg.scala 16:16]
  reg  r_269; // @[Reg.scala 16:16]
  reg  r_270; // @[Reg.scala 16:16]
  reg  r_271; // @[Reg.scala 16:16]
  reg  r_272; // @[Reg.scala 16:16]
  reg  r_273; // @[Reg.scala 16:16]
  reg  r_274; // @[Reg.scala 16:16]
  reg  r_275; // @[Reg.scala 16:16]
  reg  r_276; // @[Reg.scala 16:16]
  reg  r_277; // @[Reg.scala 16:16]
  reg  r_278; // @[Reg.scala 16:16]
  reg  r_279; // @[Reg.scala 16:16]
  reg  r_280; // @[Reg.scala 16:16]
  reg  r_281; // @[Reg.scala 16:16]
  reg  r_282; // @[Reg.scala 16:16]
  reg  r_283; // @[Reg.scala 16:16]
  reg  r_284; // @[Reg.scala 16:16]
  reg  r_285; // @[Reg.scala 16:16]
  reg  r_286; // @[Reg.scala 16:16]
  reg  r_287; // @[Reg.scala 16:16]
  reg  r_288; // @[Reg.scala 16:16]
  reg  r_289; // @[Reg.scala 16:16]
  reg  r_290; // @[Reg.scala 16:16]
  reg  r_291; // @[Reg.scala 16:16]
  reg  r_292; // @[Reg.scala 16:16]
  reg  r_293; // @[Reg.scala 16:16]
  reg  r_294; // @[Reg.scala 16:16]
  reg  r_295; // @[Reg.scala 16:16]
  reg  r_296; // @[Reg.scala 16:16]
  reg  r_297; // @[Reg.scala 16:16]
  reg  r_298; // @[Reg.scala 16:16]
  reg  r_299; // @[Reg.scala 16:16]
  reg  r_300; // @[Reg.scala 16:16]
  reg  r_301; // @[Reg.scala 16:16]
  reg  r_302; // @[Reg.scala 16:16]
  reg  r_303; // @[Reg.scala 16:16]
  reg  r_304; // @[Reg.scala 16:16]
  reg  r_305; // @[Reg.scala 16:16]
  reg  r_306; // @[Reg.scala 16:16]
  reg  r_307; // @[Reg.scala 16:16]
  reg  r_308; // @[Reg.scala 16:16]
  reg  r_309; // @[Reg.scala 16:16]
  reg  r_310; // @[Reg.scala 16:16]
  reg  r_311; // @[Reg.scala 16:16]
  reg  r_312; // @[Reg.scala 16:16]
  reg  r_313; // @[Reg.scala 16:16]
  reg  r_314; // @[Reg.scala 16:16]
  reg  r_315; // @[Reg.scala 16:16]
  reg  r_316; // @[Reg.scala 16:16]
  reg  r_317; // @[Reg.scala 16:16]
  reg  r_318; // @[Reg.scala 16:16]
  reg  r_319; // @[Reg.scala 16:16]
  reg  r_320; // @[Reg.scala 16:16]
  reg  r_321; // @[Reg.scala 16:16]
  reg  r_322; // @[Reg.scala 16:16]
  reg  r_323; // @[Reg.scala 16:16]
  reg  r_324; // @[Reg.scala 16:16]
  reg  r_325; // @[Reg.scala 16:16]
  reg  r_326; // @[Reg.scala 16:16]
  reg  r_327; // @[Reg.scala 16:16]
  reg  r_328; // @[Reg.scala 16:16]
  reg  r_329; // @[Reg.scala 16:16]
  reg  r_330; // @[Reg.scala 16:16]
  reg  r_331; // @[Reg.scala 16:16]
  reg  r_332; // @[Reg.scala 16:16]
  reg  r_333; // @[Reg.scala 16:16]
  reg  r_334; // @[Reg.scala 16:16]
  reg  r_335; // @[Reg.scala 16:16]
  reg  r_336; // @[Reg.scala 16:16]
  reg  r_337; // @[Reg.scala 16:16]
  reg  r_338; // @[Reg.scala 16:16]
  reg  r_339; // @[Reg.scala 16:16]
  reg  r_340; // @[Reg.scala 16:16]
  reg  r_341; // @[Reg.scala 16:16]
  reg  r_342; // @[Reg.scala 16:16]
  reg  r_343; // @[Reg.scala 16:16]
  reg  r_344; // @[Reg.scala 16:16]
  reg  r_345; // @[Reg.scala 16:16]
  reg  r_346; // @[Reg.scala 16:16]
  reg  r_347; // @[Reg.scala 16:16]
  reg  r_348; // @[Reg.scala 16:16]
  reg  r_349; // @[Reg.scala 16:16]
  reg  r_350; // @[Reg.scala 16:16]
  reg  r_351; // @[Reg.scala 16:16]
  reg  r_352; // @[Reg.scala 16:16]
  reg  r_353; // @[Reg.scala 16:16]
  reg  r_354; // @[Reg.scala 16:16]
  reg  r_355; // @[Reg.scala 16:16]
  reg  r_356; // @[Reg.scala 16:16]
  reg  r_357; // @[Reg.scala 16:16]
  reg  r_358; // @[Reg.scala 16:16]
  reg  r_359; // @[Reg.scala 16:16]
  reg  r_360; // @[Reg.scala 16:16]
  reg  r_361; // @[Reg.scala 16:16]
  reg  r_362; // @[Reg.scala 16:16]
  reg  r_363; // @[Reg.scala 16:16]
  reg  r_364; // @[Reg.scala 16:16]
  reg  r_365; // @[Reg.scala 16:16]
  reg  r_366; // @[Reg.scala 16:16]
  reg  r_367; // @[Reg.scala 16:16]
  reg  r_368; // @[Reg.scala 16:16]
  reg  r_369; // @[Reg.scala 16:16]
  reg  r_370; // @[Reg.scala 16:16]
  reg  r_371; // @[Reg.scala 16:16]
  reg  r_372; // @[Reg.scala 16:16]
  reg  r_373; // @[Reg.scala 16:16]
  reg  r_374; // @[Reg.scala 16:16]
  reg  r_375; // @[Reg.scala 16:16]
  reg  r_376; // @[Reg.scala 16:16]
  reg  r_377; // @[Reg.scala 16:16]
  reg  r_378; // @[Reg.scala 16:16]
  reg  r_379; // @[Reg.scala 16:16]
  reg  r_380; // @[Reg.scala 16:16]
  reg  r_381; // @[Reg.scala 16:16]
  reg  r_382; // @[Reg.scala 16:16]
  reg  r_383; // @[Reg.scala 16:16]
  reg  r_384; // @[Reg.scala 16:16]
  reg  r_385; // @[Reg.scala 16:16]
  reg  r_386; // @[Reg.scala 16:16]
  reg  r_387; // @[Reg.scala 16:16]
  reg  r_388; // @[Reg.scala 16:16]
  reg  r_389; // @[Reg.scala 16:16]
  reg  r_390; // @[Reg.scala 16:16]
  reg  r_391; // @[Reg.scala 16:16]
  reg  r_392; // @[Reg.scala 16:16]
  reg  r_393; // @[Reg.scala 16:16]
  reg  r_394; // @[Reg.scala 16:16]
  reg  r_395; // @[Reg.scala 16:16]
  reg  r_396; // @[Reg.scala 16:16]
  reg  r_397; // @[Reg.scala 16:16]
  reg  r_398; // @[Reg.scala 16:16]
  reg  r_399; // @[Reg.scala 16:16]
  reg  r_400; // @[Reg.scala 16:16]
  reg  r_401; // @[Reg.scala 16:16]
  reg  r_402; // @[Reg.scala 16:16]
  reg  r_403; // @[Reg.scala 16:16]
  reg  r_404; // @[Reg.scala 16:16]
  reg  r_405; // @[Reg.scala 16:16]
  reg  r_406; // @[Reg.scala 16:16]
  reg  r_407; // @[Reg.scala 16:16]
  reg  r_408; // @[Reg.scala 16:16]
  reg  r_409; // @[Reg.scala 16:16]
  reg  r_410; // @[Reg.scala 16:16]
  reg  r_411; // @[Reg.scala 16:16]
  reg  r_412; // @[Reg.scala 16:16]
  reg  r_413; // @[Reg.scala 16:16]
  reg  r_414; // @[Reg.scala 16:16]
  reg  r_415; // @[Reg.scala 16:16]
  reg  r_416; // @[Reg.scala 16:16]
  reg  r_417; // @[Reg.scala 16:16]
  reg  r_418; // @[Reg.scala 16:16]
  reg  r_419; // @[Reg.scala 16:16]
  reg  r_420; // @[Reg.scala 16:16]
  reg  r_421; // @[Reg.scala 16:16]
  reg  r_422; // @[Reg.scala 16:16]
  reg  r_423; // @[Reg.scala 16:16]
  reg  r_424; // @[Reg.scala 16:16]
  reg  r_425; // @[Reg.scala 16:16]
  reg  r_426; // @[Reg.scala 16:16]
  reg  r_427; // @[Reg.scala 16:16]
  reg  r_428; // @[Reg.scala 16:16]
  reg  r_429; // @[Reg.scala 16:16]
  reg  r_430; // @[Reg.scala 16:16]
  reg  r_431; // @[Reg.scala 16:16]
  reg  r_432; // @[Reg.scala 16:16]
  reg  r_433; // @[Reg.scala 16:16]
  reg  r_434; // @[Reg.scala 16:16]
  reg  r_435; // @[Reg.scala 16:16]
  reg  r_436; // @[Reg.scala 16:16]
  reg  r_437; // @[Reg.scala 16:16]
  reg  r_438; // @[Reg.scala 16:16]
  reg  r_439; // @[Reg.scala 16:16]
  reg  r_440; // @[Reg.scala 16:16]
  reg  r_441; // @[Reg.scala 16:16]
  reg  r_442; // @[Reg.scala 16:16]
  reg  r_443; // @[Reg.scala 16:16]
  reg  r_444; // @[Reg.scala 16:16]
  reg  r_445; // @[Reg.scala 16:16]
  reg  r_446; // @[Reg.scala 16:16]
  reg  r_447; // @[Reg.scala 16:16]
  reg  r_448; // @[Reg.scala 16:16]
  reg  r_449; // @[Reg.scala 16:16]
  reg  r_450; // @[Reg.scala 16:16]
  reg  r_451; // @[Reg.scala 16:16]
  reg  r_452; // @[Reg.scala 16:16]
  reg  r_453; // @[Reg.scala 16:16]
  reg  r_454; // @[Reg.scala 16:16]
  reg  r_455; // @[Reg.scala 16:16]
  reg  r_456; // @[Reg.scala 16:16]
  reg  r_457; // @[Reg.scala 16:16]
  reg  r_458; // @[Reg.scala 16:16]
  reg  r_459; // @[Reg.scala 16:16]
  reg  r_460; // @[Reg.scala 16:16]
  reg  r_461; // @[Reg.scala 16:16]
  reg  r_462; // @[Reg.scala 16:16]
  reg  r_463; // @[Reg.scala 16:16]
  reg  r_464; // @[Reg.scala 16:16]
  reg  r_465; // @[Reg.scala 16:16]
  reg  r_466; // @[Reg.scala 16:16]
  reg  r_467; // @[Reg.scala 16:16]
  reg  r_468; // @[Reg.scala 16:16]
  reg  r_469; // @[Reg.scala 16:16]
  reg  r_470; // @[Reg.scala 16:16]
  reg  r_471; // @[Reg.scala 16:16]
  reg  r_472; // @[Reg.scala 16:16]
  reg  r_473; // @[Reg.scala 16:16]
  reg  r_474; // @[Reg.scala 16:16]
  reg  r_475; // @[Reg.scala 16:16]
  reg  r_476; // @[Reg.scala 16:16]
  reg  r_477; // @[Reg.scala 16:16]
  reg  r_478; // @[Reg.scala 16:16]
  reg  r_479; // @[Reg.scala 16:16]
  reg  r_480; // @[Reg.scala 16:16]
  reg  r_481; // @[Reg.scala 16:16]
  reg  r_482; // @[Reg.scala 16:16]
  reg  r_483; // @[Reg.scala 16:16]
  reg  r_484; // @[Reg.scala 16:16]
  reg  r_485; // @[Reg.scala 16:16]
  reg  r_486; // @[Reg.scala 16:16]
  reg  r_487; // @[Reg.scala 16:16]
  reg  r_488; // @[Reg.scala 16:16]
  reg  r_489; // @[Reg.scala 16:16]
  reg  r_490; // @[Reg.scala 16:16]
  reg  r_491; // @[Reg.scala 16:16]
  reg  r_492; // @[Reg.scala 16:16]
  reg  r_493; // @[Reg.scala 16:16]
  reg  r_494; // @[Reg.scala 16:16]
  reg  r_495; // @[Reg.scala 16:16]
  reg  r_496; // @[Reg.scala 16:16]
  reg  r_497; // @[Reg.scala 16:16]
  reg  r_498; // @[Reg.scala 16:16]
  reg  r_499; // @[Reg.scala 16:16]
  reg  r_500; // @[Reg.scala 16:16]
  reg  r_501; // @[Reg.scala 16:16]
  reg  r_502; // @[Reg.scala 16:16]
  reg  r_503; // @[Reg.scala 16:16]
  reg  r_504; // @[Reg.scala 16:16]
  reg  r_505; // @[Reg.scala 16:16]
  reg  r_506; // @[Reg.scala 16:16]
  reg  r_507; // @[Reg.scala 16:16]
  reg  r_508; // @[Reg.scala 16:16]
  reg  r_509; // @[Reg.scala 16:16]
  reg  r_510; // @[Reg.scala 16:16]
  reg  r_511; // @[Reg.scala 16:16]
  reg  r_512; // @[Reg.scala 16:16]
  reg  r_513; // @[Reg.scala 16:16]
  reg  r_514; // @[Reg.scala 16:16]
  reg  r_515; // @[Reg.scala 16:16]
  reg  r_516; // @[Reg.scala 16:16]
  reg  r_517; // @[Reg.scala 16:16]
  reg  r_518; // @[Reg.scala 16:16]
  reg  r_519; // @[Reg.scala 16:16]
  reg  r_520; // @[Reg.scala 16:16]
  reg  r_521; // @[Reg.scala 16:16]
  reg  r_522; // @[Reg.scala 16:16]
  reg  r_523; // @[Reg.scala 16:16]
  reg  r_524; // @[Reg.scala 16:16]
  reg  r_525; // @[Reg.scala 16:16]
  reg  r_526; // @[Reg.scala 16:16]
  reg  r_527; // @[Reg.scala 16:16]
  reg  r_528; // @[Reg.scala 16:16]
  reg  r_529; // @[Reg.scala 16:16]
  reg  r_530; // @[Reg.scala 16:16]
  reg  r_531; // @[Reg.scala 16:16]
  reg  r_532; // @[Reg.scala 16:16]
  reg  r_533; // @[Reg.scala 16:16]
  reg  r_534; // @[Reg.scala 16:16]
  reg  r_535; // @[Reg.scala 16:16]
  reg  r_536; // @[Reg.scala 16:16]
  reg  r_537; // @[Reg.scala 16:16]
  reg  r_538; // @[Reg.scala 16:16]
  reg  r_539; // @[Reg.scala 16:16]
  reg  r_540; // @[Reg.scala 16:16]
  reg  r_541; // @[Reg.scala 16:16]
  reg  r_542; // @[Reg.scala 16:16]
  reg  r_543; // @[Reg.scala 16:16]
  reg  r_544; // @[Reg.scala 16:16]
  reg  r_545; // @[Reg.scala 16:16]
  reg  r_546; // @[Reg.scala 16:16]
  reg  r_547; // @[Reg.scala 16:16]
  reg  r_548; // @[Reg.scala 16:16]
  reg  r_549; // @[Reg.scala 16:16]
  reg  r_550; // @[Reg.scala 16:16]
  reg  r_551; // @[Reg.scala 16:16]
  reg  r_552; // @[Reg.scala 16:16]
  reg  r_553; // @[Reg.scala 16:16]
  reg  r_554; // @[Reg.scala 16:16]
  reg  r_555; // @[Reg.scala 16:16]
  reg  r_556; // @[Reg.scala 16:16]
  reg  r_557; // @[Reg.scala 16:16]
  reg  r_558; // @[Reg.scala 16:16]
  reg  r_559; // @[Reg.scala 16:16]
  reg  r_560; // @[Reg.scala 16:16]
  reg  r_561; // @[Reg.scala 16:16]
  reg  r_562; // @[Reg.scala 16:16]
  reg  r_563; // @[Reg.scala 16:16]
  reg  r_564; // @[Reg.scala 16:16]
  reg  r_565; // @[Reg.scala 16:16]
  reg  r_566; // @[Reg.scala 16:16]
  reg  r_567; // @[Reg.scala 16:16]
  reg  r_568; // @[Reg.scala 16:16]
  reg  r_569; // @[Reg.scala 16:16]
  reg  r_570; // @[Reg.scala 16:16]
  reg  r_571; // @[Reg.scala 16:16]
  reg  r_572; // @[Reg.scala 16:16]
  reg  r_573; // @[Reg.scala 16:16]
  reg  r_574; // @[Reg.scala 16:16]
  reg  r_575; // @[Reg.scala 16:16]
  reg  r_576; // @[Reg.scala 16:16]
  reg  r_577; // @[Reg.scala 16:16]
  reg  r_578; // @[Reg.scala 16:16]
  reg  r_579; // @[Reg.scala 16:16]
  reg  r_580; // @[Reg.scala 16:16]
  reg  r_581; // @[Reg.scala 16:16]
  reg  r_582; // @[Reg.scala 16:16]
  reg  r_583; // @[Reg.scala 16:16]
  reg  r_584; // @[Reg.scala 16:16]
  reg  r_585; // @[Reg.scala 16:16]
  reg  r_586; // @[Reg.scala 16:16]
  reg  r_587; // @[Reg.scala 16:16]
  reg  r_588; // @[Reg.scala 16:16]
  reg  r_589; // @[Reg.scala 16:16]
  reg  r_590; // @[Reg.scala 16:16]
  reg  r_591; // @[Reg.scala 16:16]
  reg  r_592; // @[Reg.scala 16:16]
  reg  r_593; // @[Reg.scala 16:16]
  reg  r_594; // @[Reg.scala 16:16]
  reg  r_595; // @[Reg.scala 16:16]
  reg  r_596; // @[Reg.scala 16:16]
  reg  r_597; // @[Reg.scala 16:16]
  reg  r_598; // @[Reg.scala 16:16]
  reg  r_599; // @[Reg.scala 16:16]
  reg  r_600; // @[Reg.scala 16:16]
  reg  r_601; // @[Reg.scala 16:16]
  reg  r_602; // @[Reg.scala 16:16]
  reg  r_603; // @[Reg.scala 16:16]
  reg  r_604; // @[Reg.scala 16:16]
  reg  r_605; // @[Reg.scala 16:16]
  reg  r_606; // @[Reg.scala 16:16]
  reg  r_607; // @[Reg.scala 16:16]
  reg  r_608; // @[Reg.scala 16:16]
  reg  r_609; // @[Reg.scala 16:16]
  reg  r_610; // @[Reg.scala 16:16]
  reg  r_611; // @[Reg.scala 16:16]
  reg  r_612; // @[Reg.scala 16:16]
  reg  r_613; // @[Reg.scala 16:16]
  reg  r_614; // @[Reg.scala 16:16]
  reg  r_615; // @[Reg.scala 16:16]
  reg  r_616; // @[Reg.scala 16:16]
  reg  r_617; // @[Reg.scala 16:16]
  reg  r_618; // @[Reg.scala 16:16]
  reg  r_619; // @[Reg.scala 16:16]
  reg  r_620; // @[Reg.scala 16:16]
  reg  r_621; // @[Reg.scala 16:16]
  reg  r_622; // @[Reg.scala 16:16]
  reg  r_623; // @[Reg.scala 16:16]
  reg  r_624; // @[Reg.scala 16:16]
  reg  r_625; // @[Reg.scala 16:16]
  reg  r_626; // @[Reg.scala 16:16]
  reg  r_627; // @[Reg.scala 16:16]
  reg  r_628; // @[Reg.scala 16:16]
  reg  r_629; // @[Reg.scala 16:16]
  reg  r_630; // @[Reg.scala 16:16]
  reg  r_631; // @[Reg.scala 16:16]
  reg  r_632; // @[Reg.scala 16:16]
  reg  r_633; // @[Reg.scala 16:16]
  reg  r_634; // @[Reg.scala 16:16]
  reg  r_635; // @[Reg.scala 16:16]
  reg  r_636; // @[Reg.scala 16:16]
  reg  r_637; // @[Reg.scala 16:16]
  reg  r_638; // @[Reg.scala 16:16]
  reg  r_639; // @[Reg.scala 16:16]
  reg  r_640; // @[Reg.scala 16:16]
  reg  r_641; // @[Reg.scala 16:16]
  reg  r_642; // @[Reg.scala 16:16]
  reg  r_643; // @[Reg.scala 16:16]
  reg  r_644; // @[Reg.scala 16:16]
  reg  r_645; // @[Reg.scala 16:16]
  reg  r_646; // @[Reg.scala 16:16]
  reg  r_647; // @[Reg.scala 16:16]
  reg  r_648; // @[Reg.scala 16:16]
  reg  r_649; // @[Reg.scala 16:16]
  reg  r_650; // @[Reg.scala 16:16]
  reg  r_651; // @[Reg.scala 16:16]
  reg  r_652; // @[Reg.scala 16:16]
  reg  r_653; // @[Reg.scala 16:16]
  reg  r_654; // @[Reg.scala 16:16]
  reg  r_655; // @[Reg.scala 16:16]
  reg  r_656; // @[Reg.scala 16:16]
  reg  r_657; // @[Reg.scala 16:16]
  reg  r_658; // @[Reg.scala 16:16]
  reg  r_659; // @[Reg.scala 16:16]
  reg  r_660; // @[Reg.scala 16:16]
  reg  r_661; // @[Reg.scala 16:16]
  reg  r_662; // @[Reg.scala 16:16]
  reg  r_663; // @[Reg.scala 16:16]
  reg  r_664; // @[Reg.scala 16:16]
  reg  r_665; // @[Reg.scala 16:16]
  reg  r_666; // @[Reg.scala 16:16]
  reg  r_667; // @[Reg.scala 16:16]
  reg  r_668; // @[Reg.scala 16:16]
  reg  r_669; // @[Reg.scala 16:16]
  reg  r_670; // @[Reg.scala 16:16]
  reg  r_671; // @[Reg.scala 16:16]
  reg  r_672; // @[Reg.scala 16:16]
  reg  r_673; // @[Reg.scala 16:16]
  reg  r_674; // @[Reg.scala 16:16]
  reg  r_675; // @[Reg.scala 16:16]
  reg  r_676; // @[Reg.scala 16:16]
  reg  r_677; // @[Reg.scala 16:16]
  reg  r_678; // @[Reg.scala 16:16]
  reg  r_679; // @[Reg.scala 16:16]
  reg  r_680; // @[Reg.scala 16:16]
  reg  r_681; // @[Reg.scala 16:16]
  reg  r_682; // @[Reg.scala 16:16]
  reg  r_683; // @[Reg.scala 16:16]
  reg  r_684; // @[Reg.scala 16:16]
  reg  r_685; // @[Reg.scala 16:16]
  reg  r_686; // @[Reg.scala 16:16]
  reg  r_687; // @[Reg.scala 16:16]
  reg  r_688; // @[Reg.scala 16:16]
  reg  r_689; // @[Reg.scala 16:16]
  reg  r_690; // @[Reg.scala 16:16]
  reg  r_691; // @[Reg.scala 16:16]
  reg  r_692; // @[Reg.scala 16:16]
  reg  r_693; // @[Reg.scala 16:16]
  reg  r_694; // @[Reg.scala 16:16]
  reg  r_695; // @[Reg.scala 16:16]
  reg  r_696; // @[Reg.scala 16:16]
  reg  r_697; // @[Reg.scala 16:16]
  reg  r_698; // @[Reg.scala 16:16]
  reg  r_699; // @[Reg.scala 16:16]
  reg  r_700; // @[Reg.scala 16:16]
  reg  r_701; // @[Reg.scala 16:16]
  reg  r_702; // @[Reg.scala 16:16]
  reg  r_703; // @[Reg.scala 16:16]
  reg  r_704; // @[Reg.scala 16:16]
  reg  r_705; // @[Reg.scala 16:16]
  reg  r_706; // @[Reg.scala 16:16]
  reg  r_707; // @[Reg.scala 16:16]
  reg  r_708; // @[Reg.scala 16:16]
  reg  r_709; // @[Reg.scala 16:16]
  reg  r_710; // @[Reg.scala 16:16]
  reg  r_711; // @[Reg.scala 16:16]
  reg  r_712; // @[Reg.scala 16:16]
  reg  r_713; // @[Reg.scala 16:16]
  reg  r_714; // @[Reg.scala 16:16]
  reg  r_715; // @[Reg.scala 16:16]
  reg  r_716; // @[Reg.scala 16:16]
  reg  r_717; // @[Reg.scala 16:16]
  reg  r_718; // @[Reg.scala 16:16]
  reg  r_719; // @[Reg.scala 16:16]
  reg  r_720; // @[Reg.scala 16:16]
  reg  r_721; // @[Reg.scala 16:16]
  reg  r_722; // @[Reg.scala 16:16]
  reg  r_723; // @[Reg.scala 16:16]
  reg  r_724; // @[Reg.scala 16:16]
  reg  r_725; // @[Reg.scala 16:16]
  reg  r_726; // @[Reg.scala 16:16]
  reg  r_727; // @[Reg.scala 16:16]
  reg  r_728; // @[Reg.scala 16:16]
  reg  r_729; // @[Reg.scala 16:16]
  reg  r_730; // @[Reg.scala 16:16]
  reg  r_731; // @[Reg.scala 16:16]
  reg  r_732; // @[Reg.scala 16:16]
  reg  r_733; // @[Reg.scala 16:16]
  reg  r_734; // @[Reg.scala 16:16]
  reg  r_735; // @[Reg.scala 16:16]
  reg  r_736; // @[Reg.scala 16:16]
  reg  r_737; // @[Reg.scala 16:16]
  reg  r_738; // @[Reg.scala 16:16]
  reg  r_739; // @[Reg.scala 16:16]
  reg  r_740; // @[Reg.scala 16:16]
  reg  r_741; // @[Reg.scala 16:16]
  reg  r_742; // @[Reg.scala 16:16]
  reg  r_743; // @[Reg.scala 16:16]
  reg  r_744; // @[Reg.scala 16:16]
  reg  r_745; // @[Reg.scala 16:16]
  reg  r_746; // @[Reg.scala 16:16]
  reg  r_747; // @[Reg.scala 16:16]
  reg  r_748; // @[Reg.scala 16:16]
  reg  r_749; // @[Reg.scala 16:16]
  reg  r_750; // @[Reg.scala 16:16]
  reg  r_751; // @[Reg.scala 16:16]
  reg  r_752; // @[Reg.scala 16:16]
  reg  r_753; // @[Reg.scala 16:16]
  reg  r_754; // @[Reg.scala 16:16]
  reg  r_755; // @[Reg.scala 16:16]
  reg  r_756; // @[Reg.scala 16:16]
  reg  r_757; // @[Reg.scala 16:16]
  reg  r_758; // @[Reg.scala 16:16]
  reg  r_759; // @[Reg.scala 16:16]
  reg  r_760; // @[Reg.scala 16:16]
  reg  r_761; // @[Reg.scala 16:16]
  reg  r_762; // @[Reg.scala 16:16]
  reg  r_763; // @[Reg.scala 16:16]
  reg  r_764; // @[Reg.scala 16:16]
  reg  r_765; // @[Reg.scala 16:16]
  reg  r_766; // @[Reg.scala 16:16]
  reg  r_767; // @[Reg.scala 16:16]
  reg  r_768; // @[Reg.scala 16:16]
  reg  r_769; // @[Reg.scala 16:16]
  reg  r_770; // @[Reg.scala 16:16]
  reg  r_771; // @[Reg.scala 16:16]
  reg  r_772; // @[Reg.scala 16:16]
  reg  r_773; // @[Reg.scala 16:16]
  reg  r_774; // @[Reg.scala 16:16]
  reg  r_775; // @[Reg.scala 16:16]
  reg  r_776; // @[Reg.scala 16:16]
  reg  r_777; // @[Reg.scala 16:16]
  reg  r_778; // @[Reg.scala 16:16]
  reg  r_779; // @[Reg.scala 16:16]
  reg  r_780; // @[Reg.scala 16:16]
  reg  r_781; // @[Reg.scala 16:16]
  reg  r_782; // @[Reg.scala 16:16]
  reg  r_783; // @[Reg.scala 16:16]
  reg  r_784; // @[Reg.scala 16:16]
  reg  r_785; // @[Reg.scala 16:16]
  reg  r_786; // @[Reg.scala 16:16]
  reg  r_787; // @[Reg.scala 16:16]
  reg  r_788; // @[Reg.scala 16:16]
  reg  r_789; // @[Reg.scala 16:16]
  reg  r_790; // @[Reg.scala 16:16]
  reg  r_791; // @[Reg.scala 16:16]
  reg  r_792; // @[Reg.scala 16:16]
  reg  r_793; // @[Reg.scala 16:16]
  reg  r_794; // @[Reg.scala 16:16]
  reg  r_795; // @[Reg.scala 16:16]
  reg  r_796; // @[Reg.scala 16:16]
  reg  r_797; // @[Reg.scala 16:16]
  reg  r_798; // @[Reg.scala 16:16]
  reg  r_799; // @[Reg.scala 16:16]
  reg  r_800; // @[Reg.scala 16:16]
  reg  r_801; // @[Reg.scala 16:16]
  reg  r_802; // @[Reg.scala 16:16]
  reg  r_803; // @[Reg.scala 16:16]
  reg  r_804; // @[Reg.scala 16:16]
  reg  r_805; // @[Reg.scala 16:16]
  reg  r_806; // @[Reg.scala 16:16]
  reg  r_807; // @[Reg.scala 16:16]
  reg  r_808; // @[Reg.scala 16:16]
  reg  r_809; // @[Reg.scala 16:16]
  reg  r_810; // @[Reg.scala 16:16]
  reg  r_811; // @[Reg.scala 16:16]
  reg  r_812; // @[Reg.scala 16:16]
  reg  r_813; // @[Reg.scala 16:16]
  reg  r_814; // @[Reg.scala 16:16]
  reg  r_815; // @[Reg.scala 16:16]
  reg  r_816; // @[Reg.scala 16:16]
  reg  r_817; // @[Reg.scala 16:16]
  reg  r_818; // @[Reg.scala 16:16]
  reg  r_819; // @[Reg.scala 16:16]
  reg  r_820; // @[Reg.scala 16:16]
  reg  r_821; // @[Reg.scala 16:16]
  reg  r_822; // @[Reg.scala 16:16]
  reg  r_823; // @[Reg.scala 16:16]
  reg  r_824; // @[Reg.scala 16:16]
  reg  r_825; // @[Reg.scala 16:16]
  reg  r_826; // @[Reg.scala 16:16]
  reg  r_827; // @[Reg.scala 16:16]
  reg  r_828; // @[Reg.scala 16:16]
  reg  r_829; // @[Reg.scala 16:16]
  reg  r_830; // @[Reg.scala 16:16]
  reg  r_831; // @[Reg.scala 16:16]
  reg  r_832; // @[Reg.scala 16:16]
  reg  r_833; // @[Reg.scala 16:16]
  reg  r_834; // @[Reg.scala 16:16]
  reg  r_835; // @[Reg.scala 16:16]
  reg  r_836; // @[Reg.scala 16:16]
  reg  r_837; // @[Reg.scala 16:16]
  reg  r_838; // @[Reg.scala 16:16]
  reg  r_839; // @[Reg.scala 16:16]
  reg  r_840; // @[Reg.scala 16:16]
  reg  r_841; // @[Reg.scala 16:16]
  reg  r_842; // @[Reg.scala 16:16]
  reg  r_843; // @[Reg.scala 16:16]
  reg  r_844; // @[Reg.scala 16:16]
  reg  r_845; // @[Reg.scala 16:16]
  reg  r_846; // @[Reg.scala 16:16]
  reg  r_847; // @[Reg.scala 16:16]
  reg  r_848; // @[Reg.scala 16:16]
  reg  r_849; // @[Reg.scala 16:16]
  reg  r_850; // @[Reg.scala 16:16]
  reg  r_851; // @[Reg.scala 16:16]
  reg  r_852; // @[Reg.scala 16:16]
  reg  r_853; // @[Reg.scala 16:16]
  reg  r_854; // @[Reg.scala 16:16]
  reg  r_855; // @[Reg.scala 16:16]
  reg  r_856; // @[Reg.scala 16:16]
  reg  r_857; // @[Reg.scala 16:16]
  reg  r_858; // @[Reg.scala 16:16]
  reg  r_859; // @[Reg.scala 16:16]
  reg  r_860; // @[Reg.scala 16:16]
  reg  r_861; // @[Reg.scala 16:16]
  reg  r_862; // @[Reg.scala 16:16]
  reg  r_863; // @[Reg.scala 16:16]
  reg  r_864; // @[Reg.scala 16:16]
  reg  r_865; // @[Reg.scala 16:16]
  reg  r_866; // @[Reg.scala 16:16]
  reg  r_867; // @[Reg.scala 16:16]
  reg  r_868; // @[Reg.scala 16:16]
  reg  r_869; // @[Reg.scala 16:16]
  reg  r_870; // @[Reg.scala 16:16]
  reg  r_871; // @[Reg.scala 16:16]
  reg  r_872; // @[Reg.scala 16:16]
  reg  r_873; // @[Reg.scala 16:16]
  reg  r_874; // @[Reg.scala 16:16]
  reg  r_875; // @[Reg.scala 16:16]
  reg  r_876; // @[Reg.scala 16:16]
  reg  r_877; // @[Reg.scala 16:16]
  reg  r_878; // @[Reg.scala 16:16]
  reg  r_879; // @[Reg.scala 16:16]
  reg  r_880; // @[Reg.scala 16:16]
  reg  r_881; // @[Reg.scala 16:16]
  reg  r_882; // @[Reg.scala 16:16]
  reg  r_883; // @[Reg.scala 16:16]
  reg  r_884; // @[Reg.scala 16:16]
  reg  r_885; // @[Reg.scala 16:16]
  reg  r_886; // @[Reg.scala 16:16]
  reg  r_887; // @[Reg.scala 16:16]
  reg  r_888; // @[Reg.scala 16:16]
  reg  r_889; // @[Reg.scala 16:16]
  reg  r_890; // @[Reg.scala 16:16]
  reg  r_891; // @[Reg.scala 16:16]
  reg  r_892; // @[Reg.scala 16:16]
  reg  r_893; // @[Reg.scala 16:16]
  reg  r_894; // @[Reg.scala 16:16]
  reg  r_895; // @[Reg.scala 16:16]
  reg  r_896; // @[Reg.scala 16:16]
  reg  r_897; // @[Reg.scala 16:16]
  reg  r_898; // @[Reg.scala 16:16]
  reg  r_899; // @[Reg.scala 16:16]
  reg  r_900; // @[Reg.scala 16:16]
  reg  r_901; // @[Reg.scala 16:16]
  reg  r_902; // @[Reg.scala 16:16]
  reg  r_903; // @[Reg.scala 16:16]
  reg  r_904; // @[Reg.scala 16:16]
  reg  r_905; // @[Reg.scala 16:16]
  reg  r_906; // @[Reg.scala 16:16]
  reg  r_907; // @[Reg.scala 16:16]
  reg  r_908; // @[Reg.scala 16:16]
  reg  r_909; // @[Reg.scala 16:16]
  reg  r_910; // @[Reg.scala 16:16]
  reg  r_911; // @[Reg.scala 16:16]
  reg  r_912; // @[Reg.scala 16:16]
  reg  r_913; // @[Reg.scala 16:16]
  reg  r_914; // @[Reg.scala 16:16]
  reg  r_915; // @[Reg.scala 16:16]
  reg  r_916; // @[Reg.scala 16:16]
  reg  r_917; // @[Reg.scala 16:16]
  reg  r_918; // @[Reg.scala 16:16]
  reg  r_919; // @[Reg.scala 16:16]
  reg  r_920; // @[Reg.scala 16:16]
  reg  r_921; // @[Reg.scala 16:16]
  reg  r_922; // @[Reg.scala 16:16]
  reg  r_923; // @[Reg.scala 16:16]
  reg  r_924; // @[Reg.scala 16:16]
  reg  r_925; // @[Reg.scala 16:16]
  reg  r_926; // @[Reg.scala 16:16]
  reg  r_927; // @[Reg.scala 16:16]
  reg  r_928; // @[Reg.scala 16:16]
  reg  r_929; // @[Reg.scala 16:16]
  reg  r_930; // @[Reg.scala 16:16]
  reg  r_931; // @[Reg.scala 16:16]
  reg  r_932; // @[Reg.scala 16:16]
  reg  r_933; // @[Reg.scala 16:16]
  reg  r_934; // @[Reg.scala 16:16]
  reg  r_935; // @[Reg.scala 16:16]
  reg  r_936; // @[Reg.scala 16:16]
  reg  r_937; // @[Reg.scala 16:16]
  reg  r_938; // @[Reg.scala 16:16]
  reg  r_939; // @[Reg.scala 16:16]
  reg  r_940; // @[Reg.scala 16:16]
  reg  r_941; // @[Reg.scala 16:16]
  reg  r_942; // @[Reg.scala 16:16]
  reg  r_943; // @[Reg.scala 16:16]
  reg  r_944; // @[Reg.scala 16:16]
  reg  r_945; // @[Reg.scala 16:16]
  reg  r_946; // @[Reg.scala 16:16]
  reg  r_947; // @[Reg.scala 16:16]
  reg  r_948; // @[Reg.scala 16:16]
  reg  r_949; // @[Reg.scala 16:16]
  reg  r_950; // @[Reg.scala 16:16]
  reg  r_951; // @[Reg.scala 16:16]
  reg  r_952; // @[Reg.scala 16:16]
  reg  r_953; // @[Reg.scala 16:16]
  reg  r_954; // @[Reg.scala 16:16]
  reg  r_955; // @[Reg.scala 16:16]
  reg  r_956; // @[Reg.scala 16:16]
  reg  r_957; // @[Reg.scala 16:16]
  reg  r_958; // @[Reg.scala 16:16]
  reg  r_959; // @[Reg.scala 16:16]
  reg  r_960; // @[Reg.scala 16:16]
  reg  r_961; // @[Reg.scala 16:16]
  reg  r_962; // @[Reg.scala 16:16]
  reg  r_963; // @[Reg.scala 16:16]
  reg  r_964; // @[Reg.scala 16:16]
  reg  r_965; // @[Reg.scala 16:16]
  reg  r_966; // @[Reg.scala 16:16]
  reg  r_967; // @[Reg.scala 16:16]
  reg  r_968; // @[Reg.scala 16:16]
  reg  r_969; // @[Reg.scala 16:16]
  reg  r_970; // @[Reg.scala 16:16]
  reg  r_971; // @[Reg.scala 16:16]
  reg  r_972; // @[Reg.scala 16:16]
  reg  r_973; // @[Reg.scala 16:16]
  reg  r_974; // @[Reg.scala 16:16]
  reg  r_975; // @[Reg.scala 16:16]
  reg  r_976; // @[Reg.scala 16:16]
  reg  r_977; // @[Reg.scala 16:16]
  reg  r_978; // @[Reg.scala 16:16]
  reg  r_979; // @[Reg.scala 16:16]
  reg  r_980; // @[Reg.scala 16:16]
  reg  r_981; // @[Reg.scala 16:16]
  reg  r_982; // @[Reg.scala 16:16]
  reg  r_983; // @[Reg.scala 16:16]
  reg  r_984; // @[Reg.scala 16:16]
  reg  r_985; // @[Reg.scala 16:16]
  reg  r_986; // @[Reg.scala 16:16]
  reg  r_987; // @[Reg.scala 16:16]
  reg  r_988; // @[Reg.scala 16:16]
  reg  r_989; // @[Reg.scala 16:16]
  reg  r_990; // @[Reg.scala 16:16]
  reg  r_991; // @[Reg.scala 16:16]
  reg  r_992; // @[Reg.scala 16:16]
  reg  r_993; // @[Reg.scala 16:16]
  reg  r_994; // @[Reg.scala 16:16]
  reg  r_995; // @[Reg.scala 16:16]
  reg  r_996; // @[Reg.scala 16:16]
  reg  r_997; // @[Reg.scala 16:16]
  reg  r_998; // @[Reg.scala 16:16]
  reg  r_999; // @[Reg.scala 16:16]
  reg  r_1000; // @[Reg.scala 16:16]
  reg  r_1001; // @[Reg.scala 16:16]
  reg  r_1002; // @[Reg.scala 16:16]
  reg  r_1003; // @[Reg.scala 16:16]
  reg  r_1004; // @[Reg.scala 16:16]
  reg  r_1005; // @[Reg.scala 16:16]
  reg  r_1006; // @[Reg.scala 16:16]
  reg  r_1007; // @[Reg.scala 16:16]
  reg  r_1008; // @[Reg.scala 16:16]
  reg  r_1009; // @[Reg.scala 16:16]
  reg  r_1010; // @[Reg.scala 16:16]
  reg  r_1011; // @[Reg.scala 16:16]
  reg  r_1012; // @[Reg.scala 16:16]
  reg  r_1013; // @[Reg.scala 16:16]
  reg  r_1014; // @[Reg.scala 16:16]
  reg  r_1015; // @[Reg.scala 16:16]
  reg  r_1016; // @[Reg.scala 16:16]
  reg  r_1017; // @[Reg.scala 16:16]
  reg  r_1018; // @[Reg.scala 16:16]
  reg  r_1019; // @[Reg.scala 16:16]
  reg  r_1020; // @[Reg.scala 16:16]
  reg  r_1021; // @[Reg.scala 16:16]
  reg  r_1022; // @[Reg.scala 16:16]
  reg  r_1023; // @[Reg.scala 16:16]
  reg  r_1024; // @[Reg.scala 16:16]
  reg  r_1025; // @[Reg.scala 16:16]
  reg  r_1026; // @[Reg.scala 16:16]
  reg  r_1027; // @[Reg.scala 16:16]
  reg  r_1028; // @[Reg.scala 16:16]
  reg  r_1029; // @[Reg.scala 16:16]
  reg  r_1030; // @[Reg.scala 16:16]
  reg  r_1031; // @[Reg.scala 16:16]
  reg  r_1032; // @[Reg.scala 16:16]
  reg  r_1033; // @[Reg.scala 16:16]
  reg  r_1034; // @[Reg.scala 16:16]
  reg  r_1035; // @[Reg.scala 16:16]
  reg  r_1036; // @[Reg.scala 16:16]
  reg  r_1037; // @[Reg.scala 16:16]
  reg  r_1038; // @[Reg.scala 16:16]
  reg  r_1039; // @[Reg.scala 16:16]
  reg  r_1040; // @[Reg.scala 16:16]
  reg  r_1041; // @[Reg.scala 16:16]
  reg  r_1042; // @[Reg.scala 16:16]
  reg  r_1043; // @[Reg.scala 16:16]
  reg  r_1044; // @[Reg.scala 16:16]
  reg  r_1045; // @[Reg.scala 16:16]
  reg  r_1046; // @[Reg.scala 16:16]
  reg  r_1047; // @[Reg.scala 16:16]
  reg  r_1048; // @[Reg.scala 16:16]
  reg  r_1049; // @[Reg.scala 16:16]
  reg  r_1050; // @[Reg.scala 16:16]
  reg  r_1051; // @[Reg.scala 16:16]
  reg  r_1052; // @[Reg.scala 16:16]
  reg  r_1053; // @[Reg.scala 16:16]
  reg  r_1054; // @[Reg.scala 16:16]
  reg  r_1055; // @[Reg.scala 16:16]
  reg  r_1056; // @[Reg.scala 16:16]
  reg  r_1057; // @[Reg.scala 16:16]
  reg  r_1058; // @[Reg.scala 16:16]
  reg  r_1059; // @[Reg.scala 16:16]
  reg  r_1060; // @[Reg.scala 16:16]
  reg  r_1061; // @[Reg.scala 16:16]
  reg  r_1062; // @[Reg.scala 16:16]
  reg  r_1063; // @[Reg.scala 16:16]
  reg  r_1064; // @[Reg.scala 16:16]
  reg  r_1065; // @[Reg.scala 16:16]
  reg  r_1066; // @[Reg.scala 16:16]
  reg  r_1067; // @[Reg.scala 16:16]
  reg  r_1068; // @[Reg.scala 16:16]
  reg  r_1069; // @[Reg.scala 16:16]
  reg  r_1070; // @[Reg.scala 16:16]
  reg  r_1071; // @[Reg.scala 16:16]
  reg  r_1072; // @[Reg.scala 16:16]
  reg  r_1073; // @[Reg.scala 16:16]
  reg  r_1074; // @[Reg.scala 16:16]
  reg  r_1075; // @[Reg.scala 16:16]
  reg  r_1076; // @[Reg.scala 16:16]
  reg  r_1077; // @[Reg.scala 16:16]
  reg  r_1078; // @[Reg.scala 16:16]
  reg  r_1079; // @[Reg.scala 16:16]
  reg  r_1080; // @[Reg.scala 16:16]
  reg  r_1081; // @[Reg.scala 16:16]
  reg  r_1082; // @[Reg.scala 16:16]
  reg  r_1083; // @[Reg.scala 16:16]
  reg  r_1084; // @[Reg.scala 16:16]
  reg  r_1085; // @[Reg.scala 16:16]
  reg  r_1086; // @[Reg.scala 16:16]
  reg  r_1087; // @[Reg.scala 16:16]
  reg  r_1088; // @[Reg.scala 16:16]
  reg  r_1089; // @[Reg.scala 16:16]
  reg  r_1090; // @[Reg.scala 16:16]
  reg  r_1091; // @[Reg.scala 16:16]
  reg  r_1092; // @[Reg.scala 16:16]
  reg  r_1093; // @[Reg.scala 16:16]
  reg  r_1094; // @[Reg.scala 16:16]
  reg  r_1095; // @[Reg.scala 16:16]
  reg  r_1096; // @[Reg.scala 16:16]
  reg  r_1097; // @[Reg.scala 16:16]
  reg  r_1098; // @[Reg.scala 16:16]
  reg  r_1099; // @[Reg.scala 16:16]
  reg  r_1100; // @[Reg.scala 16:16]
  reg  r_1101; // @[Reg.scala 16:16]
  reg  r_1102; // @[Reg.scala 16:16]
  reg  r_1103; // @[Reg.scala 16:16]
  reg  r_1104; // @[Reg.scala 16:16]
  reg  r_1105; // @[Reg.scala 16:16]
  reg  r_1106; // @[Reg.scala 16:16]
  reg  r_1107; // @[Reg.scala 16:16]
  reg  r_1108; // @[Reg.scala 16:16]
  reg  r_1109; // @[Reg.scala 16:16]
  reg  r_1110; // @[Reg.scala 16:16]
  reg  r_1111; // @[Reg.scala 16:16]
  reg  r_1112; // @[Reg.scala 16:16]
  reg  r_1113; // @[Reg.scala 16:16]
  reg  r_1114; // @[Reg.scala 16:16]
  reg  r_1115; // @[Reg.scala 16:16]
  reg  r_1116; // @[Reg.scala 16:16]
  reg  r_1117; // @[Reg.scala 16:16]
  reg  r_1118; // @[Reg.scala 16:16]
  reg  r_1119; // @[Reg.scala 16:16]
  reg  r_1120; // @[Reg.scala 16:16]
  reg  r_1121; // @[Reg.scala 16:16]
  reg  r_1122; // @[Reg.scala 16:16]
  reg  r_1123; // @[Reg.scala 16:16]
  reg  r_1124; // @[Reg.scala 16:16]
  reg  r_1125; // @[Reg.scala 16:16]
  reg  r_1126; // @[Reg.scala 16:16]
  reg  r_1127; // @[Reg.scala 16:16]
  reg  r_1128; // @[Reg.scala 16:16]
  reg  r_1129; // @[Reg.scala 16:16]
  reg  r_1130; // @[Reg.scala 16:16]
  reg  r_1131; // @[Reg.scala 16:16]
  reg  r_1132; // @[Reg.scala 16:16]
  reg  r_1133; // @[Reg.scala 16:16]
  reg  r_1134; // @[Reg.scala 16:16]
  reg  r_1135; // @[Reg.scala 16:16]
  reg  r_1136; // @[Reg.scala 16:16]
  reg  r_1137; // @[Reg.scala 16:16]
  reg  r_1138; // @[Reg.scala 16:16]
  reg  r_1139; // @[Reg.scala 16:16]
  reg  r_1140; // @[Reg.scala 16:16]
  reg  r_1141; // @[Reg.scala 16:16]
  reg  r_1142; // @[Reg.scala 16:16]
  reg  r_1143; // @[Reg.scala 16:16]
  reg  r_1144; // @[Reg.scala 16:16]
  reg  r_1145; // @[Reg.scala 16:16]
  reg  r_1146; // @[Reg.scala 16:16]
  reg  r_1147; // @[Reg.scala 16:16]
  reg  r_1148; // @[Reg.scala 16:16]
  reg  r_1149; // @[Reg.scala 16:16]
  reg  r_1150; // @[Reg.scala 16:16]
  reg  r_1151; // @[Reg.scala 16:16]
  reg  r_1152; // @[Reg.scala 16:16]
  reg  r_1153; // @[Reg.scala 16:16]
  reg  r_1154; // @[Reg.scala 16:16]
  reg  r_1155; // @[Reg.scala 16:16]
  reg  r_1156; // @[Reg.scala 16:16]
  reg  r_1157; // @[Reg.scala 16:16]
  reg  r_1158; // @[Reg.scala 16:16]
  reg  r_1159; // @[Reg.scala 16:16]
  reg  r_1160; // @[Reg.scala 16:16]
  reg  r_1161; // @[Reg.scala 16:16]
  reg  r_1162; // @[Reg.scala 16:16]
  reg  r_1163; // @[Reg.scala 16:16]
  reg  r_1164; // @[Reg.scala 16:16]
  reg  r_1165; // @[Reg.scala 16:16]
  reg  r_1166; // @[Reg.scala 16:16]
  reg  r_1167; // @[Reg.scala 16:16]
  reg  r_1168; // @[Reg.scala 16:16]
  reg  r_1169; // @[Reg.scala 16:16]
  reg  r_1170; // @[Reg.scala 16:16]
  reg  r_1171; // @[Reg.scala 16:16]
  reg  r_1172; // @[Reg.scala 16:16]
  reg  r_1173; // @[Reg.scala 16:16]
  reg  r_1174; // @[Reg.scala 16:16]
  reg  r_1175; // @[Reg.scala 16:16]
  reg  r_1176; // @[Reg.scala 16:16]
  reg  r_1177; // @[Reg.scala 16:16]
  reg  r_1178; // @[Reg.scala 16:16]
  reg  r_1179; // @[Reg.scala 16:16]
  reg  r_1180; // @[Reg.scala 16:16]
  reg  r_1181; // @[Reg.scala 16:16]
  reg  r_1182; // @[Reg.scala 16:16]
  reg  r_1183; // @[Reg.scala 16:16]
  reg  r_1184; // @[Reg.scala 16:16]
  reg  r_1185; // @[Reg.scala 16:16]
  reg  r_1186; // @[Reg.scala 16:16]
  reg  r_1187; // @[Reg.scala 16:16]
  reg  r_1188; // @[Reg.scala 16:16]
  reg  r_1189; // @[Reg.scala 16:16]
  reg  r_1190; // @[Reg.scala 16:16]
  reg  r_1191; // @[Reg.scala 16:16]
  reg  r_1192; // @[Reg.scala 16:16]
  reg  r_1193; // @[Reg.scala 16:16]
  reg  r_1194; // @[Reg.scala 16:16]
  reg  r_1195; // @[Reg.scala 16:16]
  reg  r_1196; // @[Reg.scala 16:16]
  reg  r_1197; // @[Reg.scala 16:16]
  reg  r_1198; // @[Reg.scala 16:16]
  reg  r_1199; // @[Reg.scala 16:16]
  reg  r_1200; // @[Reg.scala 16:16]
  reg  r_1201; // @[Reg.scala 16:16]
  reg  r_1202; // @[Reg.scala 16:16]
  reg  r_1203; // @[Reg.scala 16:16]
  reg  r_1204; // @[Reg.scala 16:16]
  reg  r_1205; // @[Reg.scala 16:16]
  reg  r_1206; // @[Reg.scala 16:16]
  reg  r_1207; // @[Reg.scala 16:16]
  reg  r_1208; // @[Reg.scala 16:16]
  reg  r_1209; // @[Reg.scala 16:16]
  reg  r_1210; // @[Reg.scala 16:16]
  reg  r_1211; // @[Reg.scala 16:16]
  reg  r_1212; // @[Reg.scala 16:16]
  reg  r_1213; // @[Reg.scala 16:16]
  reg  r_1214; // @[Reg.scala 16:16]
  reg  r_1215; // @[Reg.scala 16:16]
  reg  r_1216; // @[Reg.scala 16:16]
  reg  r_1217; // @[Reg.scala 16:16]
  reg  r_1218; // @[Reg.scala 16:16]
  reg  r_1219; // @[Reg.scala 16:16]
  reg  r_1220; // @[Reg.scala 16:16]
  reg  r_1221; // @[Reg.scala 16:16]
  reg  r_1222; // @[Reg.scala 16:16]
  reg  r_1223; // @[Reg.scala 16:16]
  reg  r_1224; // @[Reg.scala 16:16]
  reg  r_1225; // @[Reg.scala 16:16]
  reg  r_1226; // @[Reg.scala 16:16]
  reg  r_1227; // @[Reg.scala 16:16]
  reg  r_1228; // @[Reg.scala 16:16]
  reg  r_1229; // @[Reg.scala 16:16]
  reg  r_1230; // @[Reg.scala 16:16]
  reg  r_1231; // @[Reg.scala 16:16]
  reg  r_1232; // @[Reg.scala 16:16]
  reg  r_1233; // @[Reg.scala 16:16]
  reg  r_1234; // @[Reg.scala 16:16]
  reg  r_1235; // @[Reg.scala 16:16]
  reg  r_1236; // @[Reg.scala 16:16]
  reg  r_1237; // @[Reg.scala 16:16]
  reg  r_1238; // @[Reg.scala 16:16]
  reg  r_1239; // @[Reg.scala 16:16]
  reg  r_1240; // @[Reg.scala 16:16]
  reg  r_1241; // @[Reg.scala 16:16]
  reg  r_1242; // @[Reg.scala 16:16]
  reg  r_1243; // @[Reg.scala 16:16]
  reg  r_1244; // @[Reg.scala 16:16]
  reg  r_1245; // @[Reg.scala 16:16]
  reg  r_1246; // @[Reg.scala 16:16]
  reg  r_1247; // @[Reg.scala 16:16]
  reg  r_1248; // @[Reg.scala 16:16]
  reg  r_1249; // @[Reg.scala 16:16]
  reg  r_1250; // @[Reg.scala 16:16]
  reg  r_1251; // @[Reg.scala 16:16]
  reg  r_1252; // @[Reg.scala 16:16]
  reg  r_1253; // @[Reg.scala 16:16]
  reg  r_1254; // @[Reg.scala 16:16]
  reg  r_1255; // @[Reg.scala 16:16]
  reg  r_1256; // @[Reg.scala 16:16]
  reg  r_1257; // @[Reg.scala 16:16]
  reg  r_1258; // @[Reg.scala 16:16]
  reg  r_1259; // @[Reg.scala 16:16]
  reg  r_1260; // @[Reg.scala 16:16]
  reg  r_1261; // @[Reg.scala 16:16]
  reg  r_1262; // @[Reg.scala 16:16]
  reg  r_1263; // @[Reg.scala 16:16]
  reg  r_1264; // @[Reg.scala 16:16]
  reg  r_1265; // @[Reg.scala 16:16]
  reg  r_1266; // @[Reg.scala 16:16]
  reg  r_1267; // @[Reg.scala 16:16]
  reg  r_1268; // @[Reg.scala 16:16]
  reg  r_1269; // @[Reg.scala 16:16]
  reg  r_1270; // @[Reg.scala 16:16]
  reg  r_1271; // @[Reg.scala 16:16]
  reg  r_1272; // @[Reg.scala 16:16]
  reg  r_1273; // @[Reg.scala 16:16]
  reg  r_1274; // @[Reg.scala 16:16]
  reg  r_1275; // @[Reg.scala 16:16]
  reg  r_1276; // @[Reg.scala 16:16]
  reg  r_1277; // @[Reg.scala 16:16]
  reg  r_1278; // @[Reg.scala 16:16]
  reg  r_1279; // @[Reg.scala 16:16]
  reg  r_1280; // @[Reg.scala 16:16]
  reg  r_1281; // @[Reg.scala 16:16]
  reg  r_1282; // @[Reg.scala 16:16]
  reg  r_1283; // @[Reg.scala 16:16]
  reg  r_1284; // @[Reg.scala 16:16]
  reg  r_1286; // @[Reg.scala 16:16]
  reg  r_1287; // @[Reg.scala 16:16]
  reg  r_1288; // @[Reg.scala 16:16]
  reg  r_1289; // @[Reg.scala 16:16]
  reg  r_1290; // @[Reg.scala 16:16]
  reg  r_1291; // @[Reg.scala 16:16]
  reg  r_1292; // @[Reg.scala 16:16]
  reg  r_1293; // @[Reg.scala 16:16]
  reg  r_1294; // @[Reg.scala 16:16]
  reg  r_1295; // @[Reg.scala 16:16]
  reg  r_1296; // @[Reg.scala 16:16]
  reg  r_1297; // @[Reg.scala 16:16]
  reg  r_1298; // @[Reg.scala 16:16]
  reg  r_1299; // @[Reg.scala 16:16]
  reg  r_1300; // @[Reg.scala 16:16]
  reg  r_1301; // @[Reg.scala 16:16]
  reg  r_1302; // @[Reg.scala 16:16]
  reg  r_1303; // @[Reg.scala 16:16]
  reg  r_1304; // @[Reg.scala 16:16]
  reg  r_1305; // @[Reg.scala 16:16]
  reg  r_1306; // @[Reg.scala 16:16]
  reg  r_1307; // @[Reg.scala 16:16]
  reg  r_1308; // @[Reg.scala 16:16]
  reg  r_1309; // @[Reg.scala 16:16]
  reg  r_1310; // @[Reg.scala 16:16]
  reg  r_1311; // @[Reg.scala 16:16]
  reg  r_1312; // @[Reg.scala 16:16]
  reg  r_1313; // @[Reg.scala 16:16]
  reg  r_1314; // @[Reg.scala 16:16]
  reg  r_1315; // @[Reg.scala 16:16]
  reg  r_1316; // @[Reg.scala 16:16]
  reg  r_1317; // @[Reg.scala 16:16]
  reg  r_1318; // @[Reg.scala 16:16]
  reg  r_1319; // @[Reg.scala 16:16]
  reg  r_1320; // @[Reg.scala 16:16]
  reg  r_1321; // @[Reg.scala 16:16]
  reg  r_1322; // @[Reg.scala 16:16]
  reg  r_1323; // @[Reg.scala 16:16]
  reg  r_1324; // @[Reg.scala 16:16]
  reg  r_1325; // @[Reg.scala 16:16]
  reg  r_1326; // @[Reg.scala 16:16]
  reg  r_1327; // @[Reg.scala 16:16]
  reg  r_1328; // @[Reg.scala 16:16]
  reg  r_1329; // @[Reg.scala 16:16]
  reg  r_1330; // @[Reg.scala 16:16]
  reg  r_1331; // @[Reg.scala 16:16]
  reg  r_1332; // @[Reg.scala 16:16]
  reg  r_1333; // @[Reg.scala 16:16]
  reg  r_1334; // @[Reg.scala 16:16]
  reg  r_1335; // @[Reg.scala 16:16]
  reg  r_1336; // @[Reg.scala 16:16]
  reg  r_1337; // @[Reg.scala 16:16]
  reg  r_1338; // @[Reg.scala 16:16]
  reg  r_1339; // @[Reg.scala 16:16]
  reg  r_1340; // @[Reg.scala 16:16]
  reg  r_1341; // @[Reg.scala 16:16]
  reg  r_1342; // @[Reg.scala 16:16]
  reg  r_1343; // @[Reg.scala 16:16]
  reg  r_1344; // @[Reg.scala 16:16]
  reg  r_1345; // @[Reg.scala 16:16]
  reg  r_1346; // @[Reg.scala 16:16]
  reg  r_1347; // @[Reg.scala 16:16]
  reg  r_1349; // @[Reg.scala 16:16]
  reg  r_1350; // @[Reg.scala 16:16]
  reg  r_1351; // @[Reg.scala 16:16]
  reg  r_1352; // @[Reg.scala 16:16]
  reg  r_1353; // @[Reg.scala 16:16]
  reg  r_1354; // @[Reg.scala 16:16]
  reg  r_1355; // @[Reg.scala 16:16]
  reg  r_1356; // @[Reg.scala 16:16]
  reg  r_1357; // @[Reg.scala 16:16]
  reg  r_1358; // @[Reg.scala 16:16]
  reg  r_1359; // @[Reg.scala 16:16]
  reg  r_1360; // @[Reg.scala 16:16]
  reg  r_1361; // @[Reg.scala 16:16]
  reg  r_1362; // @[Reg.scala 16:16]
  reg  r_1363; // @[Reg.scala 16:16]
  reg  r_1364; // @[Reg.scala 16:16]
  reg  r_1365; // @[Reg.scala 16:16]
  reg  r_1366; // @[Reg.scala 16:16]
  reg  r_1367; // @[Reg.scala 16:16]
  reg  r_1368; // @[Reg.scala 16:16]
  reg  r_1369; // @[Reg.scala 16:16]
  reg  r_1370; // @[Reg.scala 16:16]
  reg  r_1371; // @[Reg.scala 16:16]
  reg  r_1372; // @[Reg.scala 16:16]
  reg  r_1373; // @[Reg.scala 16:16]
  reg  r_1374; // @[Reg.scala 16:16]
  reg  r_1375; // @[Reg.scala 16:16]
  reg  r_1376; // @[Reg.scala 16:16]
  reg  r_1377; // @[Reg.scala 16:16]
  reg  r_1378; // @[Reg.scala 16:16]
  reg  r_1379; // @[Reg.scala 16:16]
  reg  r_1380; // @[Reg.scala 16:16]
  reg  r_1381; // @[Reg.scala 16:16]
  reg  r_1382; // @[Reg.scala 16:16]
  reg  r_1383; // @[Reg.scala 16:16]
  reg  r_1384; // @[Reg.scala 16:16]
  reg  r_1385; // @[Reg.scala 16:16]
  reg  r_1386; // @[Reg.scala 16:16]
  reg  r_1387; // @[Reg.scala 16:16]
  reg  r_1388; // @[Reg.scala 16:16]
  reg  r_1389; // @[Reg.scala 16:16]
  reg  r_1390; // @[Reg.scala 16:16]
  reg  r_1391; // @[Reg.scala 16:16]
  reg  r_1392; // @[Reg.scala 16:16]
  reg  r_1393; // @[Reg.scala 16:16]
  reg  r_1394; // @[Reg.scala 16:16]
  reg  r_1395; // @[Reg.scala 16:16]
  reg  r_1396; // @[Reg.scala 16:16]
  reg  r_1397; // @[Reg.scala 16:16]
  reg  r_1398; // @[Reg.scala 16:16]
  reg  r_1399; // @[Reg.scala 16:16]
  reg  r_1400; // @[Reg.scala 16:16]
  reg  r_1401; // @[Reg.scala 16:16]
  reg  r_1402; // @[Reg.scala 16:16]
  reg  r_1403; // @[Reg.scala 16:16]
  reg  r_1404; // @[Reg.scala 16:16]
  reg  r_1405; // @[Reg.scala 16:16]
  reg  r_1406; // @[Reg.scala 16:16]
  reg  r_1407; // @[Reg.scala 16:16]
  reg  r_1408; // @[Reg.scala 16:16]
  reg  r_1410; // @[Reg.scala 16:16]
  reg  r_1411; // @[Reg.scala 16:16]
  reg  r_1412; // @[Reg.scala 16:16]
  reg  r_1413; // @[Reg.scala 16:16]
  reg  r_1414; // @[Reg.scala 16:16]
  reg  r_1415; // @[Reg.scala 16:16]
  reg  r_1416; // @[Reg.scala 16:16]
  reg  r_1417; // @[Reg.scala 16:16]
  reg  r_1418; // @[Reg.scala 16:16]
  reg  r_1419; // @[Reg.scala 16:16]
  reg  r_1420; // @[Reg.scala 16:16]
  reg  r_1421; // @[Reg.scala 16:16]
  reg  r_1422; // @[Reg.scala 16:16]
  reg  r_1423; // @[Reg.scala 16:16]
  reg  r_1424; // @[Reg.scala 16:16]
  reg  r_1425; // @[Reg.scala 16:16]
  reg  r_1426; // @[Reg.scala 16:16]
  reg  r_1427; // @[Reg.scala 16:16]
  reg  r_1428; // @[Reg.scala 16:16]
  reg  r_1429; // @[Reg.scala 16:16]
  reg  r_1430; // @[Reg.scala 16:16]
  reg  r_1431; // @[Reg.scala 16:16]
  reg  r_1432; // @[Reg.scala 16:16]
  reg  r_1433; // @[Reg.scala 16:16]
  reg  r_1434; // @[Reg.scala 16:16]
  reg  r_1435; // @[Reg.scala 16:16]
  reg  r_1436; // @[Reg.scala 16:16]
  reg  r_1437; // @[Reg.scala 16:16]
  reg  r_1438; // @[Reg.scala 16:16]
  reg  r_1439; // @[Reg.scala 16:16]
  reg  r_1440; // @[Reg.scala 16:16]
  reg  r_1441; // @[Reg.scala 16:16]
  reg  r_1442; // @[Reg.scala 16:16]
  reg  r_1443; // @[Reg.scala 16:16]
  reg  r_1444; // @[Reg.scala 16:16]
  reg  r_1445; // @[Reg.scala 16:16]
  reg  r_1446; // @[Reg.scala 16:16]
  reg  r_1447; // @[Reg.scala 16:16]
  reg  r_1448; // @[Reg.scala 16:16]
  reg  r_1449; // @[Reg.scala 16:16]
  reg  r_1450; // @[Reg.scala 16:16]
  reg  r_1451; // @[Reg.scala 16:16]
  reg  r_1452; // @[Reg.scala 16:16]
  reg  r_1453; // @[Reg.scala 16:16]
  reg  r_1454; // @[Reg.scala 16:16]
  reg  r_1455; // @[Reg.scala 16:16]
  reg  r_1456; // @[Reg.scala 16:16]
  reg  r_1457; // @[Reg.scala 16:16]
  reg  r_1458; // @[Reg.scala 16:16]
  reg  r_1459; // @[Reg.scala 16:16]
  reg  r_1460; // @[Reg.scala 16:16]
  reg  r_1461; // @[Reg.scala 16:16]
  reg  r_1462; // @[Reg.scala 16:16]
  reg  r_1463; // @[Reg.scala 16:16]
  reg  r_1464; // @[Reg.scala 16:16]
  reg  r_1465; // @[Reg.scala 16:16]
  reg  r_1466; // @[Reg.scala 16:16]
  reg  r_1467; // @[Reg.scala 16:16]
  reg  r_1469; // @[Reg.scala 16:16]
  reg  r_1470; // @[Reg.scala 16:16]
  reg  r_1471; // @[Reg.scala 16:16]
  reg  r_1472; // @[Reg.scala 16:16]
  reg  r_1473; // @[Reg.scala 16:16]
  reg  r_1474; // @[Reg.scala 16:16]
  reg  r_1475; // @[Reg.scala 16:16]
  reg  r_1476; // @[Reg.scala 16:16]
  reg  r_1477; // @[Reg.scala 16:16]
  reg  r_1478; // @[Reg.scala 16:16]
  reg  r_1479; // @[Reg.scala 16:16]
  reg  r_1480; // @[Reg.scala 16:16]
  reg  r_1481; // @[Reg.scala 16:16]
  reg  r_1482; // @[Reg.scala 16:16]
  reg  r_1483; // @[Reg.scala 16:16]
  reg  r_1484; // @[Reg.scala 16:16]
  reg  r_1485; // @[Reg.scala 16:16]
  reg  r_1486; // @[Reg.scala 16:16]
  reg  r_1487; // @[Reg.scala 16:16]
  reg  r_1488; // @[Reg.scala 16:16]
  reg  r_1489; // @[Reg.scala 16:16]
  reg  r_1490; // @[Reg.scala 16:16]
  reg  r_1491; // @[Reg.scala 16:16]
  reg  r_1492; // @[Reg.scala 16:16]
  reg  r_1493; // @[Reg.scala 16:16]
  reg  r_1494; // @[Reg.scala 16:16]
  reg  r_1495; // @[Reg.scala 16:16]
  reg  r_1496; // @[Reg.scala 16:16]
  reg  r_1497; // @[Reg.scala 16:16]
  reg  r_1498; // @[Reg.scala 16:16]
  reg  r_1499; // @[Reg.scala 16:16]
  reg  r_1500; // @[Reg.scala 16:16]
  reg  r_1501; // @[Reg.scala 16:16]
  reg  r_1502; // @[Reg.scala 16:16]
  reg  r_1503; // @[Reg.scala 16:16]
  reg  r_1504; // @[Reg.scala 16:16]
  reg  r_1505; // @[Reg.scala 16:16]
  reg  r_1506; // @[Reg.scala 16:16]
  reg  r_1507; // @[Reg.scala 16:16]
  reg  r_1508; // @[Reg.scala 16:16]
  reg  r_1509; // @[Reg.scala 16:16]
  reg  r_1510; // @[Reg.scala 16:16]
  reg  r_1511; // @[Reg.scala 16:16]
  reg  r_1512; // @[Reg.scala 16:16]
  reg  r_1513; // @[Reg.scala 16:16]
  reg  r_1514; // @[Reg.scala 16:16]
  reg  r_1515; // @[Reg.scala 16:16]
  reg  r_1516; // @[Reg.scala 16:16]
  reg  r_1517; // @[Reg.scala 16:16]
  reg  r_1518; // @[Reg.scala 16:16]
  reg  r_1519; // @[Reg.scala 16:16]
  reg  r_1520; // @[Reg.scala 16:16]
  reg  r_1521; // @[Reg.scala 16:16]
  reg  r_1522; // @[Reg.scala 16:16]
  reg  r_1523; // @[Reg.scala 16:16]
  reg  r_1524; // @[Reg.scala 16:16]
  reg  r_1526; // @[Reg.scala 16:16]
  reg  r_1527; // @[Reg.scala 16:16]
  reg  r_1528; // @[Reg.scala 16:16]
  reg  r_1529; // @[Reg.scala 16:16]
  reg  r_1530; // @[Reg.scala 16:16]
  reg  r_1531; // @[Reg.scala 16:16]
  reg  r_1532; // @[Reg.scala 16:16]
  reg  r_1533; // @[Reg.scala 16:16]
  reg  r_1534; // @[Reg.scala 16:16]
  reg  r_1535; // @[Reg.scala 16:16]
  reg  r_1536; // @[Reg.scala 16:16]
  reg  r_1537; // @[Reg.scala 16:16]
  reg  r_1538; // @[Reg.scala 16:16]
  reg  r_1539; // @[Reg.scala 16:16]
  reg  r_1540; // @[Reg.scala 16:16]
  reg  r_1541; // @[Reg.scala 16:16]
  reg  r_1542; // @[Reg.scala 16:16]
  reg  r_1543; // @[Reg.scala 16:16]
  reg  r_1544; // @[Reg.scala 16:16]
  reg  r_1545; // @[Reg.scala 16:16]
  reg  r_1546; // @[Reg.scala 16:16]
  reg  r_1547; // @[Reg.scala 16:16]
  reg  r_1548; // @[Reg.scala 16:16]
  reg  r_1549; // @[Reg.scala 16:16]
  reg  r_1550; // @[Reg.scala 16:16]
  reg  r_1551; // @[Reg.scala 16:16]
  reg  r_1552; // @[Reg.scala 16:16]
  reg  r_1553; // @[Reg.scala 16:16]
  reg  r_1554; // @[Reg.scala 16:16]
  reg  r_1555; // @[Reg.scala 16:16]
  reg  r_1556; // @[Reg.scala 16:16]
  reg  r_1557; // @[Reg.scala 16:16]
  reg  r_1558; // @[Reg.scala 16:16]
  reg  r_1559; // @[Reg.scala 16:16]
  reg  r_1560; // @[Reg.scala 16:16]
  reg  r_1561; // @[Reg.scala 16:16]
  reg  r_1562; // @[Reg.scala 16:16]
  reg  r_1563; // @[Reg.scala 16:16]
  reg  r_1564; // @[Reg.scala 16:16]
  reg  r_1565; // @[Reg.scala 16:16]
  reg  r_1566; // @[Reg.scala 16:16]
  reg  r_1567; // @[Reg.scala 16:16]
  reg  r_1568; // @[Reg.scala 16:16]
  reg  r_1569; // @[Reg.scala 16:16]
  reg  r_1570; // @[Reg.scala 16:16]
  reg  r_1571; // @[Reg.scala 16:16]
  reg  r_1572; // @[Reg.scala 16:16]
  reg  r_1573; // @[Reg.scala 16:16]
  reg  r_1574; // @[Reg.scala 16:16]
  reg  r_1575; // @[Reg.scala 16:16]
  reg  r_1576; // @[Reg.scala 16:16]
  reg  r_1577; // @[Reg.scala 16:16]
  reg  r_1578; // @[Reg.scala 16:16]
  reg  r_1579; // @[Reg.scala 16:16]
  reg  r_1581; // @[Reg.scala 16:16]
  reg  r_1582; // @[Reg.scala 16:16]
  reg  r_1583; // @[Reg.scala 16:16]
  reg  r_1584; // @[Reg.scala 16:16]
  reg  r_1585; // @[Reg.scala 16:16]
  reg  r_1586; // @[Reg.scala 16:16]
  reg  r_1587; // @[Reg.scala 16:16]
  reg  r_1588; // @[Reg.scala 16:16]
  reg  r_1589; // @[Reg.scala 16:16]
  reg  r_1590; // @[Reg.scala 16:16]
  reg  r_1591; // @[Reg.scala 16:16]
  reg  r_1592; // @[Reg.scala 16:16]
  reg  r_1593; // @[Reg.scala 16:16]
  reg  r_1594; // @[Reg.scala 16:16]
  reg  r_1595; // @[Reg.scala 16:16]
  reg  r_1596; // @[Reg.scala 16:16]
  reg  r_1597; // @[Reg.scala 16:16]
  reg  r_1598; // @[Reg.scala 16:16]
  reg  r_1599; // @[Reg.scala 16:16]
  reg  r_1600; // @[Reg.scala 16:16]
  reg  r_1601; // @[Reg.scala 16:16]
  reg  r_1602; // @[Reg.scala 16:16]
  reg  r_1603; // @[Reg.scala 16:16]
  reg  r_1604; // @[Reg.scala 16:16]
  reg  r_1605; // @[Reg.scala 16:16]
  reg  r_1606; // @[Reg.scala 16:16]
  reg  r_1607; // @[Reg.scala 16:16]
  reg  r_1608; // @[Reg.scala 16:16]
  reg  r_1609; // @[Reg.scala 16:16]
  reg  r_1610; // @[Reg.scala 16:16]
  reg  r_1611; // @[Reg.scala 16:16]
  reg  r_1612; // @[Reg.scala 16:16]
  reg  r_1613; // @[Reg.scala 16:16]
  reg  r_1614; // @[Reg.scala 16:16]
  reg  r_1615; // @[Reg.scala 16:16]
  reg  r_1616; // @[Reg.scala 16:16]
  reg  r_1617; // @[Reg.scala 16:16]
  reg  r_1618; // @[Reg.scala 16:16]
  reg  r_1619; // @[Reg.scala 16:16]
  reg  r_1620; // @[Reg.scala 16:16]
  reg  r_1621; // @[Reg.scala 16:16]
  reg  r_1622; // @[Reg.scala 16:16]
  reg  r_1623; // @[Reg.scala 16:16]
  reg  r_1624; // @[Reg.scala 16:16]
  reg  r_1625; // @[Reg.scala 16:16]
  reg  r_1626; // @[Reg.scala 16:16]
  reg  r_1627; // @[Reg.scala 16:16]
  reg  r_1628; // @[Reg.scala 16:16]
  reg  r_1629; // @[Reg.scala 16:16]
  reg  r_1630; // @[Reg.scala 16:16]
  reg  r_1631; // @[Reg.scala 16:16]
  reg  r_1632; // @[Reg.scala 16:16]
  reg  r_1634; // @[Reg.scala 16:16]
  reg  r_1635; // @[Reg.scala 16:16]
  reg  r_1636; // @[Reg.scala 16:16]
  reg  r_1637; // @[Reg.scala 16:16]
  reg  r_1638; // @[Reg.scala 16:16]
  reg  r_1639; // @[Reg.scala 16:16]
  reg  r_1640; // @[Reg.scala 16:16]
  reg  r_1641; // @[Reg.scala 16:16]
  reg  r_1642; // @[Reg.scala 16:16]
  reg  r_1643; // @[Reg.scala 16:16]
  reg  r_1644; // @[Reg.scala 16:16]
  reg  r_1645; // @[Reg.scala 16:16]
  reg  r_1646; // @[Reg.scala 16:16]
  reg  r_1647; // @[Reg.scala 16:16]
  reg  r_1648; // @[Reg.scala 16:16]
  reg  r_1649; // @[Reg.scala 16:16]
  reg  r_1650; // @[Reg.scala 16:16]
  reg  r_1651; // @[Reg.scala 16:16]
  reg  r_1652; // @[Reg.scala 16:16]
  reg  r_1653; // @[Reg.scala 16:16]
  reg  r_1654; // @[Reg.scala 16:16]
  reg  r_1655; // @[Reg.scala 16:16]
  reg  r_1656; // @[Reg.scala 16:16]
  reg  r_1657; // @[Reg.scala 16:16]
  reg  r_1658; // @[Reg.scala 16:16]
  reg  r_1659; // @[Reg.scala 16:16]
  reg  r_1660; // @[Reg.scala 16:16]
  reg  r_1661; // @[Reg.scala 16:16]
  reg  r_1662; // @[Reg.scala 16:16]
  reg  r_1663; // @[Reg.scala 16:16]
  reg  r_1664; // @[Reg.scala 16:16]
  reg  r_1665; // @[Reg.scala 16:16]
  reg  r_1666; // @[Reg.scala 16:16]
  reg  r_1667; // @[Reg.scala 16:16]
  reg  r_1668; // @[Reg.scala 16:16]
  reg  r_1669; // @[Reg.scala 16:16]
  reg  r_1670; // @[Reg.scala 16:16]
  reg  r_1671; // @[Reg.scala 16:16]
  reg  r_1672; // @[Reg.scala 16:16]
  reg  r_1673; // @[Reg.scala 16:16]
  reg  r_1674; // @[Reg.scala 16:16]
  reg  r_1675; // @[Reg.scala 16:16]
  reg  r_1676; // @[Reg.scala 16:16]
  reg  r_1677; // @[Reg.scala 16:16]
  reg  r_1678; // @[Reg.scala 16:16]
  reg  r_1679; // @[Reg.scala 16:16]
  reg  r_1680; // @[Reg.scala 16:16]
  reg  r_1681; // @[Reg.scala 16:16]
  reg  r_1682; // @[Reg.scala 16:16]
  reg  r_1683; // @[Reg.scala 16:16]
  reg  r_1685; // @[Reg.scala 16:16]
  reg  r_1686; // @[Reg.scala 16:16]
  reg  r_1687; // @[Reg.scala 16:16]
  reg  r_1688; // @[Reg.scala 16:16]
  reg  r_1689; // @[Reg.scala 16:16]
  reg  r_1690; // @[Reg.scala 16:16]
  reg  r_1691; // @[Reg.scala 16:16]
  reg  r_1692; // @[Reg.scala 16:16]
  reg  r_1693; // @[Reg.scala 16:16]
  reg  r_1694; // @[Reg.scala 16:16]
  reg  r_1695; // @[Reg.scala 16:16]
  reg  r_1696; // @[Reg.scala 16:16]
  reg  r_1697; // @[Reg.scala 16:16]
  reg  r_1698; // @[Reg.scala 16:16]
  reg  r_1699; // @[Reg.scala 16:16]
  reg  r_1700; // @[Reg.scala 16:16]
  reg  r_1701; // @[Reg.scala 16:16]
  reg  r_1702; // @[Reg.scala 16:16]
  reg  r_1703; // @[Reg.scala 16:16]
  reg  r_1704; // @[Reg.scala 16:16]
  reg  r_1705; // @[Reg.scala 16:16]
  reg  r_1706; // @[Reg.scala 16:16]
  reg  r_1707; // @[Reg.scala 16:16]
  reg  r_1708; // @[Reg.scala 16:16]
  reg  r_1709; // @[Reg.scala 16:16]
  reg  r_1710; // @[Reg.scala 16:16]
  reg  r_1711; // @[Reg.scala 16:16]
  reg  r_1712; // @[Reg.scala 16:16]
  reg  r_1713; // @[Reg.scala 16:16]
  reg  r_1714; // @[Reg.scala 16:16]
  reg  r_1715; // @[Reg.scala 16:16]
  reg  r_1716; // @[Reg.scala 16:16]
  reg  r_1717; // @[Reg.scala 16:16]
  reg  r_1718; // @[Reg.scala 16:16]
  reg  r_1719; // @[Reg.scala 16:16]
  reg  r_1720; // @[Reg.scala 16:16]
  reg  r_1721; // @[Reg.scala 16:16]
  reg  r_1722; // @[Reg.scala 16:16]
  reg  r_1723; // @[Reg.scala 16:16]
  reg  r_1724; // @[Reg.scala 16:16]
  reg  r_1725; // @[Reg.scala 16:16]
  reg  r_1726; // @[Reg.scala 16:16]
  reg  r_1727; // @[Reg.scala 16:16]
  reg  r_1728; // @[Reg.scala 16:16]
  reg  r_1729; // @[Reg.scala 16:16]
  reg  r_1730; // @[Reg.scala 16:16]
  reg  r_1731; // @[Reg.scala 16:16]
  reg  r_1732; // @[Reg.scala 16:16]
  reg  r_1734; // @[Reg.scala 16:16]
  reg  r_1735; // @[Reg.scala 16:16]
  reg  r_1736; // @[Reg.scala 16:16]
  reg  r_1737; // @[Reg.scala 16:16]
  reg  r_1738; // @[Reg.scala 16:16]
  reg  r_1739; // @[Reg.scala 16:16]
  reg  r_1740; // @[Reg.scala 16:16]
  reg  r_1741; // @[Reg.scala 16:16]
  reg  r_1742; // @[Reg.scala 16:16]
  reg  r_1743; // @[Reg.scala 16:16]
  reg  r_1744; // @[Reg.scala 16:16]
  reg  r_1745; // @[Reg.scala 16:16]
  reg  r_1746; // @[Reg.scala 16:16]
  reg  r_1747; // @[Reg.scala 16:16]
  reg  r_1748; // @[Reg.scala 16:16]
  reg  r_1749; // @[Reg.scala 16:16]
  reg  r_1750; // @[Reg.scala 16:16]
  reg  r_1751; // @[Reg.scala 16:16]
  reg  r_1752; // @[Reg.scala 16:16]
  reg  r_1753; // @[Reg.scala 16:16]
  reg  r_1754; // @[Reg.scala 16:16]
  reg  r_1755; // @[Reg.scala 16:16]
  reg  r_1756; // @[Reg.scala 16:16]
  reg  r_1757; // @[Reg.scala 16:16]
  reg  r_1758; // @[Reg.scala 16:16]
  reg  r_1759; // @[Reg.scala 16:16]
  reg  r_1760; // @[Reg.scala 16:16]
  reg  r_1761; // @[Reg.scala 16:16]
  reg  r_1762; // @[Reg.scala 16:16]
  reg  r_1763; // @[Reg.scala 16:16]
  reg  r_1764; // @[Reg.scala 16:16]
  reg  r_1765; // @[Reg.scala 16:16]
  reg  r_1766; // @[Reg.scala 16:16]
  reg  r_1767; // @[Reg.scala 16:16]
  reg  r_1768; // @[Reg.scala 16:16]
  reg  r_1769; // @[Reg.scala 16:16]
  reg  r_1770; // @[Reg.scala 16:16]
  reg  r_1771; // @[Reg.scala 16:16]
  reg  r_1772; // @[Reg.scala 16:16]
  reg  r_1773; // @[Reg.scala 16:16]
  reg  r_1774; // @[Reg.scala 16:16]
  reg  r_1775; // @[Reg.scala 16:16]
  reg  r_1776; // @[Reg.scala 16:16]
  reg  r_1777; // @[Reg.scala 16:16]
  reg  r_1778; // @[Reg.scala 16:16]
  reg  r_1779; // @[Reg.scala 16:16]
  reg  r_1781; // @[Reg.scala 16:16]
  reg  r_1782; // @[Reg.scala 16:16]
  reg  r_1783; // @[Reg.scala 16:16]
  reg  r_1784; // @[Reg.scala 16:16]
  reg  r_1785; // @[Reg.scala 16:16]
  reg  r_1786; // @[Reg.scala 16:16]
  reg  r_1787; // @[Reg.scala 16:16]
  reg  r_1788; // @[Reg.scala 16:16]
  reg  r_1789; // @[Reg.scala 16:16]
  reg  r_1790; // @[Reg.scala 16:16]
  reg  r_1791; // @[Reg.scala 16:16]
  reg  r_1792; // @[Reg.scala 16:16]
  reg  r_1793; // @[Reg.scala 16:16]
  reg  r_1794; // @[Reg.scala 16:16]
  reg  r_1795; // @[Reg.scala 16:16]
  reg  r_1796; // @[Reg.scala 16:16]
  reg  r_1797; // @[Reg.scala 16:16]
  reg  r_1798; // @[Reg.scala 16:16]
  reg  r_1799; // @[Reg.scala 16:16]
  reg  r_1800; // @[Reg.scala 16:16]
  reg  r_1801; // @[Reg.scala 16:16]
  reg  r_1802; // @[Reg.scala 16:16]
  reg  r_1803; // @[Reg.scala 16:16]
  reg  r_1804; // @[Reg.scala 16:16]
  reg  r_1805; // @[Reg.scala 16:16]
  reg  r_1806; // @[Reg.scala 16:16]
  reg  r_1807; // @[Reg.scala 16:16]
  reg  r_1808; // @[Reg.scala 16:16]
  reg  r_1809; // @[Reg.scala 16:16]
  reg  r_1810; // @[Reg.scala 16:16]
  reg  r_1811; // @[Reg.scala 16:16]
  reg  r_1812; // @[Reg.scala 16:16]
  reg  r_1813; // @[Reg.scala 16:16]
  reg  r_1814; // @[Reg.scala 16:16]
  reg  r_1815; // @[Reg.scala 16:16]
  reg  r_1816; // @[Reg.scala 16:16]
  reg  r_1817; // @[Reg.scala 16:16]
  reg  r_1818; // @[Reg.scala 16:16]
  reg  r_1819; // @[Reg.scala 16:16]
  reg  r_1820; // @[Reg.scala 16:16]
  reg  r_1821; // @[Reg.scala 16:16]
  reg  r_1822; // @[Reg.scala 16:16]
  reg  r_1823; // @[Reg.scala 16:16]
  reg  r_1824; // @[Reg.scala 16:16]
  reg  r_1826; // @[Reg.scala 16:16]
  reg  r_1827; // @[Reg.scala 16:16]
  reg  r_1828; // @[Reg.scala 16:16]
  reg  r_1829; // @[Reg.scala 16:16]
  reg  r_1830; // @[Reg.scala 16:16]
  reg  r_1831; // @[Reg.scala 16:16]
  reg  r_1832; // @[Reg.scala 16:16]
  reg  r_1833; // @[Reg.scala 16:16]
  reg  r_1834; // @[Reg.scala 16:16]
  reg  r_1835; // @[Reg.scala 16:16]
  reg  r_1836; // @[Reg.scala 16:16]
  reg  r_1837; // @[Reg.scala 16:16]
  reg  r_1838; // @[Reg.scala 16:16]
  reg  r_1839; // @[Reg.scala 16:16]
  reg  r_1840; // @[Reg.scala 16:16]
  reg  r_1841; // @[Reg.scala 16:16]
  reg  r_1842; // @[Reg.scala 16:16]
  reg  r_1843; // @[Reg.scala 16:16]
  reg  r_1844; // @[Reg.scala 16:16]
  reg  r_1845; // @[Reg.scala 16:16]
  reg  r_1846; // @[Reg.scala 16:16]
  reg  r_1847; // @[Reg.scala 16:16]
  reg  r_1848; // @[Reg.scala 16:16]
  reg  r_1849; // @[Reg.scala 16:16]
  reg  r_1850; // @[Reg.scala 16:16]
  reg  r_1851; // @[Reg.scala 16:16]
  reg  r_1852; // @[Reg.scala 16:16]
  reg  r_1853; // @[Reg.scala 16:16]
  reg  r_1854; // @[Reg.scala 16:16]
  reg  r_1855; // @[Reg.scala 16:16]
  reg  r_1856; // @[Reg.scala 16:16]
  reg  r_1857; // @[Reg.scala 16:16]
  reg  r_1858; // @[Reg.scala 16:16]
  reg  r_1859; // @[Reg.scala 16:16]
  reg  r_1860; // @[Reg.scala 16:16]
  reg  r_1861; // @[Reg.scala 16:16]
  reg  r_1862; // @[Reg.scala 16:16]
  reg  r_1863; // @[Reg.scala 16:16]
  reg  r_1864; // @[Reg.scala 16:16]
  reg  r_1865; // @[Reg.scala 16:16]
  reg  r_1866; // @[Reg.scala 16:16]
  reg  r_1867; // @[Reg.scala 16:16]
  reg  r_1869; // @[Reg.scala 16:16]
  reg  r_1870; // @[Reg.scala 16:16]
  reg  r_1871; // @[Reg.scala 16:16]
  reg  r_1872; // @[Reg.scala 16:16]
  reg  r_1873; // @[Reg.scala 16:16]
  reg  r_1874; // @[Reg.scala 16:16]
  reg  r_1875; // @[Reg.scala 16:16]
  reg  r_1876; // @[Reg.scala 16:16]
  reg  r_1877; // @[Reg.scala 16:16]
  reg  r_1878; // @[Reg.scala 16:16]
  reg  r_1879; // @[Reg.scala 16:16]
  reg  r_1880; // @[Reg.scala 16:16]
  reg  r_1881; // @[Reg.scala 16:16]
  reg  r_1882; // @[Reg.scala 16:16]
  reg  r_1883; // @[Reg.scala 16:16]
  reg  r_1884; // @[Reg.scala 16:16]
  reg  r_1885; // @[Reg.scala 16:16]
  reg  r_1886; // @[Reg.scala 16:16]
  reg  r_1887; // @[Reg.scala 16:16]
  reg  r_1888; // @[Reg.scala 16:16]
  reg  r_1889; // @[Reg.scala 16:16]
  reg  r_1890; // @[Reg.scala 16:16]
  reg  r_1891; // @[Reg.scala 16:16]
  reg  r_1892; // @[Reg.scala 16:16]
  reg  r_1893; // @[Reg.scala 16:16]
  reg  r_1894; // @[Reg.scala 16:16]
  reg  r_1895; // @[Reg.scala 16:16]
  reg  r_1896; // @[Reg.scala 16:16]
  reg  r_1897; // @[Reg.scala 16:16]
  reg  r_1898; // @[Reg.scala 16:16]
  reg  r_1899; // @[Reg.scala 16:16]
  reg  r_1900; // @[Reg.scala 16:16]
  reg  r_1901; // @[Reg.scala 16:16]
  reg  r_1902; // @[Reg.scala 16:16]
  reg  r_1903; // @[Reg.scala 16:16]
  reg  r_1904; // @[Reg.scala 16:16]
  reg  r_1905; // @[Reg.scala 16:16]
  reg  r_1906; // @[Reg.scala 16:16]
  reg  r_1907; // @[Reg.scala 16:16]
  reg  r_1908; // @[Reg.scala 16:16]
  reg  r_1910; // @[Reg.scala 16:16]
  reg  r_1911; // @[Reg.scala 16:16]
  reg  r_1912; // @[Reg.scala 16:16]
  reg  r_1913; // @[Reg.scala 16:16]
  reg  r_1914; // @[Reg.scala 16:16]
  reg  r_1915; // @[Reg.scala 16:16]
  reg  r_1916; // @[Reg.scala 16:16]
  reg  r_1917; // @[Reg.scala 16:16]
  reg  r_1918; // @[Reg.scala 16:16]
  reg  r_1919; // @[Reg.scala 16:16]
  reg  r_1920; // @[Reg.scala 16:16]
  reg  r_1921; // @[Reg.scala 16:16]
  reg  r_1922; // @[Reg.scala 16:16]
  reg  r_1923; // @[Reg.scala 16:16]
  reg  r_1924; // @[Reg.scala 16:16]
  reg  r_1925; // @[Reg.scala 16:16]
  reg  r_1926; // @[Reg.scala 16:16]
  reg  r_1927; // @[Reg.scala 16:16]
  reg  r_1928; // @[Reg.scala 16:16]
  reg  r_1929; // @[Reg.scala 16:16]
  reg  r_1930; // @[Reg.scala 16:16]
  reg  r_1931; // @[Reg.scala 16:16]
  reg  r_1932; // @[Reg.scala 16:16]
  reg  r_1933; // @[Reg.scala 16:16]
  reg  r_1934; // @[Reg.scala 16:16]
  reg  r_1935; // @[Reg.scala 16:16]
  reg  r_1936; // @[Reg.scala 16:16]
  reg  r_1937; // @[Reg.scala 16:16]
  reg  r_1938; // @[Reg.scala 16:16]
  reg  r_1939; // @[Reg.scala 16:16]
  reg  r_1940; // @[Reg.scala 16:16]
  reg  r_1941; // @[Reg.scala 16:16]
  reg  r_1942; // @[Reg.scala 16:16]
  reg  r_1943; // @[Reg.scala 16:16]
  reg  r_1944; // @[Reg.scala 16:16]
  reg  r_1945; // @[Reg.scala 16:16]
  reg  r_1946; // @[Reg.scala 16:16]
  reg  r_1947; // @[Reg.scala 16:16]
  reg  r_1949; // @[Reg.scala 16:16]
  reg  r_1950; // @[Reg.scala 16:16]
  reg  r_1951; // @[Reg.scala 16:16]
  reg  r_1952; // @[Reg.scala 16:16]
  reg  r_1953; // @[Reg.scala 16:16]
  reg  r_1954; // @[Reg.scala 16:16]
  reg  r_1955; // @[Reg.scala 16:16]
  reg  r_1956; // @[Reg.scala 16:16]
  reg  r_1957; // @[Reg.scala 16:16]
  reg  r_1958; // @[Reg.scala 16:16]
  reg  r_1959; // @[Reg.scala 16:16]
  reg  r_1960; // @[Reg.scala 16:16]
  reg  r_1961; // @[Reg.scala 16:16]
  reg  r_1962; // @[Reg.scala 16:16]
  reg  r_1963; // @[Reg.scala 16:16]
  reg  r_1964; // @[Reg.scala 16:16]
  reg  r_1965; // @[Reg.scala 16:16]
  reg  r_1966; // @[Reg.scala 16:16]
  reg  r_1967; // @[Reg.scala 16:16]
  reg  r_1968; // @[Reg.scala 16:16]
  reg  r_1969; // @[Reg.scala 16:16]
  reg  r_1970; // @[Reg.scala 16:16]
  reg  r_1971; // @[Reg.scala 16:16]
  reg  r_1972; // @[Reg.scala 16:16]
  reg  r_1973; // @[Reg.scala 16:16]
  reg  r_1974; // @[Reg.scala 16:16]
  reg  r_1975; // @[Reg.scala 16:16]
  reg  r_1976; // @[Reg.scala 16:16]
  reg  r_1977; // @[Reg.scala 16:16]
  reg  r_1978; // @[Reg.scala 16:16]
  reg  r_1979; // @[Reg.scala 16:16]
  reg  r_1980; // @[Reg.scala 16:16]
  reg  r_1981; // @[Reg.scala 16:16]
  reg  r_1982; // @[Reg.scala 16:16]
  reg  r_1983; // @[Reg.scala 16:16]
  reg  r_1984; // @[Reg.scala 16:16]
  reg  r_1986; // @[Reg.scala 16:16]
  reg  r_1987; // @[Reg.scala 16:16]
  reg  r_1988; // @[Reg.scala 16:16]
  reg  r_1989; // @[Reg.scala 16:16]
  reg  r_1990; // @[Reg.scala 16:16]
  reg  r_1991; // @[Reg.scala 16:16]
  reg  r_1992; // @[Reg.scala 16:16]
  reg  r_1993; // @[Reg.scala 16:16]
  reg  r_1994; // @[Reg.scala 16:16]
  reg  r_1995; // @[Reg.scala 16:16]
  reg  r_1996; // @[Reg.scala 16:16]
  reg  r_1997; // @[Reg.scala 16:16]
  reg  r_1998; // @[Reg.scala 16:16]
  reg  r_1999; // @[Reg.scala 16:16]
  reg  r_2000; // @[Reg.scala 16:16]
  reg  r_2001; // @[Reg.scala 16:16]
  reg  r_2002; // @[Reg.scala 16:16]
  reg  r_2003; // @[Reg.scala 16:16]
  reg  r_2004; // @[Reg.scala 16:16]
  reg  r_2005; // @[Reg.scala 16:16]
  reg  r_2006; // @[Reg.scala 16:16]
  reg  r_2007; // @[Reg.scala 16:16]
  reg  r_2008; // @[Reg.scala 16:16]
  reg  r_2009; // @[Reg.scala 16:16]
  reg  r_2010; // @[Reg.scala 16:16]
  reg  r_2011; // @[Reg.scala 16:16]
  reg  r_2012; // @[Reg.scala 16:16]
  reg  r_2013; // @[Reg.scala 16:16]
  reg  r_2014; // @[Reg.scala 16:16]
  reg  r_2015; // @[Reg.scala 16:16]
  reg  r_2016; // @[Reg.scala 16:16]
  reg  r_2017; // @[Reg.scala 16:16]
  reg  r_2018; // @[Reg.scala 16:16]
  reg  r_2019; // @[Reg.scala 16:16]
  reg  r_2021; // @[Reg.scala 16:16]
  reg  r_2022; // @[Reg.scala 16:16]
  reg  r_2023; // @[Reg.scala 16:16]
  reg  r_2024; // @[Reg.scala 16:16]
  reg  r_2025; // @[Reg.scala 16:16]
  reg  r_2026; // @[Reg.scala 16:16]
  reg  r_2027; // @[Reg.scala 16:16]
  reg  r_2028; // @[Reg.scala 16:16]
  reg  r_2029; // @[Reg.scala 16:16]
  reg  r_2030; // @[Reg.scala 16:16]
  reg  r_2031; // @[Reg.scala 16:16]
  reg  r_2032; // @[Reg.scala 16:16]
  reg  r_2033; // @[Reg.scala 16:16]
  reg  r_2034; // @[Reg.scala 16:16]
  reg  r_2035; // @[Reg.scala 16:16]
  reg  r_2036; // @[Reg.scala 16:16]
  reg  r_2037; // @[Reg.scala 16:16]
  reg  r_2038; // @[Reg.scala 16:16]
  reg  r_2039; // @[Reg.scala 16:16]
  reg  r_2040; // @[Reg.scala 16:16]
  reg  r_2041; // @[Reg.scala 16:16]
  reg  r_2042; // @[Reg.scala 16:16]
  reg  r_2043; // @[Reg.scala 16:16]
  reg  r_2044; // @[Reg.scala 16:16]
  reg  r_2045; // @[Reg.scala 16:16]
  reg  r_2046; // @[Reg.scala 16:16]
  reg  r_2047; // @[Reg.scala 16:16]
  reg  r_2048; // @[Reg.scala 16:16]
  reg  r_2049; // @[Reg.scala 16:16]
  reg  r_2050; // @[Reg.scala 16:16]
  reg  r_2051; // @[Reg.scala 16:16]
  reg  r_2052; // @[Reg.scala 16:16]
  reg  r_2054; // @[Reg.scala 16:16]
  reg  r_2055; // @[Reg.scala 16:16]
  reg  r_2056; // @[Reg.scala 16:16]
  reg  r_2057; // @[Reg.scala 16:16]
  reg  r_2058; // @[Reg.scala 16:16]
  reg  r_2059; // @[Reg.scala 16:16]
  reg  r_2060; // @[Reg.scala 16:16]
  reg  r_2061; // @[Reg.scala 16:16]
  reg  r_2062; // @[Reg.scala 16:16]
  reg  r_2063; // @[Reg.scala 16:16]
  reg  r_2064; // @[Reg.scala 16:16]
  reg  r_2065; // @[Reg.scala 16:16]
  reg  r_2066; // @[Reg.scala 16:16]
  reg  r_2067; // @[Reg.scala 16:16]
  reg  r_2068; // @[Reg.scala 16:16]
  reg  r_2069; // @[Reg.scala 16:16]
  reg  r_2070; // @[Reg.scala 16:16]
  reg  r_2071; // @[Reg.scala 16:16]
  reg  r_2072; // @[Reg.scala 16:16]
  reg  r_2073; // @[Reg.scala 16:16]
  reg  r_2074; // @[Reg.scala 16:16]
  reg  r_2075; // @[Reg.scala 16:16]
  reg  r_2076; // @[Reg.scala 16:16]
  reg  r_2077; // @[Reg.scala 16:16]
  reg  r_2078; // @[Reg.scala 16:16]
  reg  r_2079; // @[Reg.scala 16:16]
  reg  r_2080; // @[Reg.scala 16:16]
  reg  r_2081; // @[Reg.scala 16:16]
  reg  r_2082; // @[Reg.scala 16:16]
  reg  r_2083; // @[Reg.scala 16:16]
  reg  r_2085; // @[Reg.scala 16:16]
  reg  r_2086; // @[Reg.scala 16:16]
  reg  r_2087; // @[Reg.scala 16:16]
  reg  r_2088; // @[Reg.scala 16:16]
  reg  r_2089; // @[Reg.scala 16:16]
  reg  r_2090; // @[Reg.scala 16:16]
  reg  r_2091; // @[Reg.scala 16:16]
  reg  r_2092; // @[Reg.scala 16:16]
  reg  r_2093; // @[Reg.scala 16:16]
  reg  r_2094; // @[Reg.scala 16:16]
  reg  r_2095; // @[Reg.scala 16:16]
  reg  r_2096; // @[Reg.scala 16:16]
  reg  r_2097; // @[Reg.scala 16:16]
  reg  r_2098; // @[Reg.scala 16:16]
  reg  r_2099; // @[Reg.scala 16:16]
  reg  r_2100; // @[Reg.scala 16:16]
  reg  r_2101; // @[Reg.scala 16:16]
  reg  r_2102; // @[Reg.scala 16:16]
  reg  r_2103; // @[Reg.scala 16:16]
  reg  r_2104; // @[Reg.scala 16:16]
  reg  r_2105; // @[Reg.scala 16:16]
  reg  r_2106; // @[Reg.scala 16:16]
  reg  r_2107; // @[Reg.scala 16:16]
  reg  r_2108; // @[Reg.scala 16:16]
  reg  r_2109; // @[Reg.scala 16:16]
  reg  r_2110; // @[Reg.scala 16:16]
  reg  r_2111; // @[Reg.scala 16:16]
  reg  r_2112; // @[Reg.scala 16:16]
  reg  r_2114; // @[Reg.scala 16:16]
  reg  r_2115; // @[Reg.scala 16:16]
  reg  r_2116; // @[Reg.scala 16:16]
  reg  r_2117; // @[Reg.scala 16:16]
  reg  r_2118; // @[Reg.scala 16:16]
  reg  r_2119; // @[Reg.scala 16:16]
  reg  r_2120; // @[Reg.scala 16:16]
  reg  r_2121; // @[Reg.scala 16:16]
  reg  r_2122; // @[Reg.scala 16:16]
  reg  r_2123; // @[Reg.scala 16:16]
  reg  r_2124; // @[Reg.scala 16:16]
  reg  r_2125; // @[Reg.scala 16:16]
  reg  r_2126; // @[Reg.scala 16:16]
  reg  r_2127; // @[Reg.scala 16:16]
  reg  r_2128; // @[Reg.scala 16:16]
  reg  r_2129; // @[Reg.scala 16:16]
  reg  r_2130; // @[Reg.scala 16:16]
  reg  r_2131; // @[Reg.scala 16:16]
  reg  r_2132; // @[Reg.scala 16:16]
  reg  r_2133; // @[Reg.scala 16:16]
  reg  r_2134; // @[Reg.scala 16:16]
  reg  r_2135; // @[Reg.scala 16:16]
  reg  r_2136; // @[Reg.scala 16:16]
  reg  r_2137; // @[Reg.scala 16:16]
  reg  r_2138; // @[Reg.scala 16:16]
  reg  r_2139; // @[Reg.scala 16:16]
  reg  r_2141; // @[Reg.scala 16:16]
  reg  r_2142; // @[Reg.scala 16:16]
  reg  r_2143; // @[Reg.scala 16:16]
  reg  r_2144; // @[Reg.scala 16:16]
  reg  r_2145; // @[Reg.scala 16:16]
  reg  r_2146; // @[Reg.scala 16:16]
  reg  r_2147; // @[Reg.scala 16:16]
  reg  r_2148; // @[Reg.scala 16:16]
  reg  r_2149; // @[Reg.scala 16:16]
  reg  r_2150; // @[Reg.scala 16:16]
  reg  r_2151; // @[Reg.scala 16:16]
  reg  r_2152; // @[Reg.scala 16:16]
  reg  r_2153; // @[Reg.scala 16:16]
  reg  r_2154; // @[Reg.scala 16:16]
  reg  r_2155; // @[Reg.scala 16:16]
  reg  r_2156; // @[Reg.scala 16:16]
  reg  r_2157; // @[Reg.scala 16:16]
  reg  r_2158; // @[Reg.scala 16:16]
  reg  r_2159; // @[Reg.scala 16:16]
  reg  r_2160; // @[Reg.scala 16:16]
  reg  r_2161; // @[Reg.scala 16:16]
  reg  r_2162; // @[Reg.scala 16:16]
  reg  r_2163; // @[Reg.scala 16:16]
  reg  r_2164; // @[Reg.scala 16:16]
  reg  r_2166; // @[Reg.scala 16:16]
  reg  r_2167; // @[Reg.scala 16:16]
  reg  r_2168; // @[Reg.scala 16:16]
  reg  r_2169; // @[Reg.scala 16:16]
  reg  r_2170; // @[Reg.scala 16:16]
  reg  r_2171; // @[Reg.scala 16:16]
  reg  r_2172; // @[Reg.scala 16:16]
  reg  r_2173; // @[Reg.scala 16:16]
  reg  r_2174; // @[Reg.scala 16:16]
  reg  r_2175; // @[Reg.scala 16:16]
  reg  r_2176; // @[Reg.scala 16:16]
  reg  r_2177; // @[Reg.scala 16:16]
  reg  r_2178; // @[Reg.scala 16:16]
  reg  r_2179; // @[Reg.scala 16:16]
  reg  r_2180; // @[Reg.scala 16:16]
  reg  r_2181; // @[Reg.scala 16:16]
  reg  r_2182; // @[Reg.scala 16:16]
  reg  r_2183; // @[Reg.scala 16:16]
  reg  r_2184; // @[Reg.scala 16:16]
  reg  r_2185; // @[Reg.scala 16:16]
  reg  r_2186; // @[Reg.scala 16:16]
  reg  r_2187; // @[Reg.scala 16:16]
  reg  r_2189; // @[Reg.scala 16:16]
  reg  r_2190; // @[Reg.scala 16:16]
  reg  r_2191; // @[Reg.scala 16:16]
  reg  r_2192; // @[Reg.scala 16:16]
  reg  r_2193; // @[Reg.scala 16:16]
  reg  r_2194; // @[Reg.scala 16:16]
  reg  r_2195; // @[Reg.scala 16:16]
  reg  r_2196; // @[Reg.scala 16:16]
  reg  r_2197; // @[Reg.scala 16:16]
  reg  r_2198; // @[Reg.scala 16:16]
  reg  r_2199; // @[Reg.scala 16:16]
  reg  r_2200; // @[Reg.scala 16:16]
  reg  r_2201; // @[Reg.scala 16:16]
  reg  r_2202; // @[Reg.scala 16:16]
  reg  r_2203; // @[Reg.scala 16:16]
  reg  r_2204; // @[Reg.scala 16:16]
  reg  r_2205; // @[Reg.scala 16:16]
  reg  r_2206; // @[Reg.scala 16:16]
  reg  r_2207; // @[Reg.scala 16:16]
  reg  r_2208; // @[Reg.scala 16:16]
  reg  r_2210; // @[Reg.scala 16:16]
  reg  r_2211; // @[Reg.scala 16:16]
  reg  r_2212; // @[Reg.scala 16:16]
  reg  r_2213; // @[Reg.scala 16:16]
  reg  r_2214; // @[Reg.scala 16:16]
  reg  r_2215; // @[Reg.scala 16:16]
  reg  r_2216; // @[Reg.scala 16:16]
  reg  r_2217; // @[Reg.scala 16:16]
  reg  r_2218; // @[Reg.scala 16:16]
  reg  r_2219; // @[Reg.scala 16:16]
  reg  r_2220; // @[Reg.scala 16:16]
  reg  r_2221; // @[Reg.scala 16:16]
  reg  r_2222; // @[Reg.scala 16:16]
  reg  r_2223; // @[Reg.scala 16:16]
  reg  r_2224; // @[Reg.scala 16:16]
  reg  r_2225; // @[Reg.scala 16:16]
  reg  r_2226; // @[Reg.scala 16:16]
  reg  r_2227; // @[Reg.scala 16:16]
  reg  r_2229; // @[Reg.scala 16:16]
  reg  r_2230; // @[Reg.scala 16:16]
  reg  r_2231; // @[Reg.scala 16:16]
  reg  r_2232; // @[Reg.scala 16:16]
  reg  r_2233; // @[Reg.scala 16:16]
  reg  r_2234; // @[Reg.scala 16:16]
  reg  r_2235; // @[Reg.scala 16:16]
  reg  r_2236; // @[Reg.scala 16:16]
  reg  r_2237; // @[Reg.scala 16:16]
  reg  r_2238; // @[Reg.scala 16:16]
  reg  r_2239; // @[Reg.scala 16:16]
  reg  r_2240; // @[Reg.scala 16:16]
  reg  r_2241; // @[Reg.scala 16:16]
  reg  r_2242; // @[Reg.scala 16:16]
  reg  r_2243; // @[Reg.scala 16:16]
  reg  r_2244; // @[Reg.scala 16:16]
  reg  r_2246; // @[Reg.scala 16:16]
  reg  r_2247; // @[Reg.scala 16:16]
  reg  r_2248; // @[Reg.scala 16:16]
  reg  r_2249; // @[Reg.scala 16:16]
  reg  r_2250; // @[Reg.scala 16:16]
  reg  r_2251; // @[Reg.scala 16:16]
  reg  r_2252; // @[Reg.scala 16:16]
  reg  r_2253; // @[Reg.scala 16:16]
  reg  r_2254; // @[Reg.scala 16:16]
  reg  r_2255; // @[Reg.scala 16:16]
  reg  r_2256; // @[Reg.scala 16:16]
  reg  r_2257; // @[Reg.scala 16:16]
  reg  r_2258; // @[Reg.scala 16:16]
  reg  r_2259; // @[Reg.scala 16:16]
  reg  r_2261; // @[Reg.scala 16:16]
  reg  r_2262; // @[Reg.scala 16:16]
  reg  r_2263; // @[Reg.scala 16:16]
  reg  r_2264; // @[Reg.scala 16:16]
  reg  r_2265; // @[Reg.scala 16:16]
  reg  r_2266; // @[Reg.scala 16:16]
  reg  r_2267; // @[Reg.scala 16:16]
  reg  r_2268; // @[Reg.scala 16:16]
  reg  r_2269; // @[Reg.scala 16:16]
  reg  r_2270; // @[Reg.scala 16:16]
  reg  r_2271; // @[Reg.scala 16:16]
  reg  r_2272; // @[Reg.scala 16:16]
  reg  r_2274; // @[Reg.scala 16:16]
  reg  r_2275; // @[Reg.scala 16:16]
  reg  r_2276; // @[Reg.scala 16:16]
  reg  r_2277; // @[Reg.scala 16:16]
  reg  r_2278; // @[Reg.scala 16:16]
  reg  r_2279; // @[Reg.scala 16:16]
  reg  r_2280; // @[Reg.scala 16:16]
  reg  r_2281; // @[Reg.scala 16:16]
  reg  r_2282; // @[Reg.scala 16:16]
  reg  r_2283; // @[Reg.scala 16:16]
  reg  r_2285; // @[Reg.scala 16:16]
  reg  r_2286; // @[Reg.scala 16:16]
  reg  r_2287; // @[Reg.scala 16:16]
  reg  r_2288; // @[Reg.scala 16:16]
  reg  r_2289; // @[Reg.scala 16:16]
  reg  r_2290; // @[Reg.scala 16:16]
  reg  r_2291; // @[Reg.scala 16:16]
  reg  r_2292; // @[Reg.scala 16:16]
  reg  r_2294; // @[Reg.scala 16:16]
  reg  r_2295; // @[Reg.scala 16:16]
  reg  r_2296; // @[Reg.scala 16:16]
  reg  r_2297; // @[Reg.scala 16:16]
  reg  r_2298; // @[Reg.scala 16:16]
  reg  r_2299; // @[Reg.scala 16:16]
  reg  r_2301; // @[Reg.scala 16:16]
  reg  r_2302; // @[Reg.scala 16:16]
  reg  r_2303; // @[Reg.scala 16:16]
  reg  r_2304; // @[Reg.scala 16:16]
  reg  r_2306; // @[Reg.scala 16:16]
  reg  r_2307; // @[Reg.scala 16:16]
  wire  c_4_78 = m_912_io_cout; // @[MUL.scala 253:22]
  wire  c_4_79 = m_917_io_cout; // @[MUL.scala 253:22]
  wire  c_4_127 = m_1217_io_cout; // @[MUL.scala 253:22]
  wire  c_1_220 = m_1352_io_cout; // @[MUL.scala 253:22]
  wire  c_1_221 = m_1354_io_cout; // @[MUL.scala 253:22]
  wire  c_1_222 = m_1356_io_cout; // @[MUL.scala 253:22]
  wire  c_1_223 = m_1358_io_cout; // @[MUL.scala 253:22]
  wire  c_4_128 = m_1492_io_cout; // @[MUL.scala 253:22]
  wire  c_4_129 = m_1497_io_cout; // @[MUL.scala 253:22]
  wire  c_4_130 = m_1502_io_cout; // @[MUL.scala 253:22]
  wire  c_4_131 = m_1507_io_cout; // @[MUL.scala 253:22]
  wire  c_4_132 = m_1512_io_cout; // @[MUL.scala 253:22]
  wire  c_4_133 = m_1517_io_cout; // @[MUL.scala 253:22]
  wire  c_4_134 = m_1522_io_cout; // @[MUL.scala 253:22]
  wire  c_4_135 = m_1527_io_cout; // @[MUL.scala 253:22]
  wire  c_4_136 = m_1532_io_cout; // @[MUL.scala 253:22]
  wire  c_4_137 = m_1537_io_cout; // @[MUL.scala 253:22]
  wire  c_1_306 = m_1666_io_cout; // @[MUL.scala 253:22]
  wire  c_1_307 = m_1668_io_cout; // @[MUL.scala 253:22]
  wire  c_1_308 = m_1670_io_cout; // @[MUL.scala 253:22]
  wire  c_1_309 = m_1672_io_cout; // @[MUL.scala 253:22]
  wire  c_1_310 = m_1674_io_cout; // @[MUL.scala 253:22]
  wire  c_1_311 = m_1676_io_cout; // @[MUL.scala 253:22]
  wire  c_1_312 = m_1678_io_cout; // @[MUL.scala 253:22]
  wire  c_1_313 = m_1680_io_cout; // @[MUL.scala 253:22]
  wire  s_0_366 = m_1706_io_s; // @[MUL.scala 252:21]
  wire  c_0_366 = m_1706_io_cout; // @[MUL.scala 253:22]
  wire  s_0_367 = m_1707_io_s; // @[MUL.scala 252:21]
  wire  c_0_367 = m_1707_io_cout; // @[MUL.scala 253:22]
  wire  s_0_368 = m_1708_io_s; // @[MUL.scala 252:21]
  wire  c_0_368 = m_1708_io_cout; // @[MUL.scala 253:22]
  wire  s_0_369 = m_1709_io_s; // @[MUL.scala 252:21]
  wire  c_0_369 = m_1709_io_cout; // @[MUL.scala 253:22]
  wire  s_0_370 = m_1710_io_s; // @[MUL.scala 252:21]
  wire  c_0_370 = m_1710_io_cout; // @[MUL.scala 253:22]
  wire  s_0_371 = m_1711_io_s; // @[MUL.scala 252:21]
  wire  c_0_371 = m_1711_io_cout; // @[MUL.scala 253:22]
  wire  s_0_372 = m_1712_io_s; // @[MUL.scala 252:21]
  wire  c_0_372 = m_1712_io_cout; // @[MUL.scala 253:22]
  wire  s_0_373 = m_1713_io_s; // @[MUL.scala 252:21]
  wire  c_0_373 = m_1713_io_cout; // @[MUL.scala 253:22]
  wire  s_0_374 = m_1714_io_s; // @[MUL.scala 252:21]
  wire  c_0_374 = m_1714_io_cout; // @[MUL.scala 253:22]
  wire  s_0_375 = m_1715_io_s; // @[MUL.scala 252:21]
  wire  c_0_375 = m_1715_io_cout; // @[MUL.scala 253:22]
  wire  s_0_376 = m_1716_io_s; // @[MUL.scala 252:21]
  wire  c_0_376 = m_1716_io_cout; // @[MUL.scala 253:22]
  wire  s_0_377 = m_1717_io_s; // @[MUL.scala 252:21]
  wire  c_0_377 = m_1717_io_cout; // @[MUL.scala 253:22]
  wire  s_0_378 = m_1718_io_s; // @[MUL.scala 252:21]
  wire  c_0_378 = m_1718_io_cout; // @[MUL.scala 253:22]
  wire  s_0_379 = m_1719_io_s; // @[MUL.scala 252:21]
  wire  c_0_379 = m_1719_io_cout; // @[MUL.scala 253:22]
  wire  s_0_380 = m_1720_io_s; // @[MUL.scala 252:21]
  wire  c_0_380 = m_1720_io_cout; // @[MUL.scala 253:22]
  wire  s_0_381 = m_1722_io_s; // @[MUL.scala 252:21]
  wire  c_0_381 = m_1722_io_cout; // @[MUL.scala 253:22]
  wire  s_0_382 = m_1724_io_s; // @[MUL.scala 252:21]
  wire  c_0_382 = m_1724_io_cout; // @[MUL.scala 253:22]
  wire  s_0_383 = m_1726_io_s; // @[MUL.scala 252:21]
  wire  c_0_383 = m_1726_io_cout; // @[MUL.scala 253:22]
  wire  s_0_384 = m_1728_io_s; // @[MUL.scala 252:21]
  wire  c_0_384 = m_1728_io_cout; // @[MUL.scala 253:22]
  wire  s_0_385 = m_1730_io_s; // @[MUL.scala 252:21]
  wire  c_0_385 = m_1730_io_cout; // @[MUL.scala 253:22]
  wire  s_2_314 = m_1731_io_s; // @[MUL.scala 252:21]
  wire  c_1_314 = m_1731_io_cout; // @[MUL.scala 253:22]
  wire  s_0_386 = m_1732_io_s; // @[MUL.scala 252:21]
  wire  c_0_386 = m_1732_io_cout; // @[MUL.scala 253:22]
  wire  s_2_315 = m_1733_io_s; // @[MUL.scala 252:21]
  wire  c_1_315 = m_1733_io_cout; // @[MUL.scala 253:22]
  wire  s_0_387 = m_1734_io_s; // @[MUL.scala 252:21]
  wire  c_0_387 = m_1734_io_cout; // @[MUL.scala 253:22]
  wire  s_2_316 = m_1735_io_s; // @[MUL.scala 252:21]
  wire  c_1_316 = m_1735_io_cout; // @[MUL.scala 253:22]
  wire  s_0_388 = m_1736_io_s; // @[MUL.scala 252:21]
  wire  c_0_388 = m_1736_io_cout; // @[MUL.scala 253:22]
  wire  s_2_317 = m_1737_io_s; // @[MUL.scala 252:21]
  wire  c_1_317 = m_1737_io_cout; // @[MUL.scala 253:22]
  wire  s_0_389 = m_1738_io_s; // @[MUL.scala 252:21]
  wire  c_0_389 = m_1738_io_cout; // @[MUL.scala 253:22]
  wire  s_2_318 = m_1739_io_s; // @[MUL.scala 252:21]
  wire  c_1_318 = m_1739_io_cout; // @[MUL.scala 253:22]
  wire  s_0_390 = m_1740_io_s; // @[MUL.scala 252:21]
  wire  c_0_390 = m_1740_io_cout; // @[MUL.scala 253:22]
  wire  s_2_319 = m_1741_io_s; // @[MUL.scala 252:21]
  wire  c_1_319 = m_1741_io_cout; // @[MUL.scala 253:22]
  wire  s_0_391 = m_1742_io_s; // @[MUL.scala 252:21]
  wire  c_0_391 = m_1742_io_cout; // @[MUL.scala 253:22]
  wire  s_2_320 = m_1743_io_s; // @[MUL.scala 252:21]
  wire  c_1_320 = m_1743_io_cout; // @[MUL.scala 253:22]
  wire  s_0_392 = m_1744_io_s; // @[MUL.scala 252:21]
  wire  c_0_392 = m_1744_io_cout; // @[MUL.scala 253:22]
  wire  s_2_321 = m_1745_io_s; // @[MUL.scala 252:21]
  wire  c_1_321 = m_1745_io_cout; // @[MUL.scala 253:22]
  wire  s_0_393 = m_1746_io_s; // @[MUL.scala 252:21]
  wire  c_0_393 = m_1746_io_cout; // @[MUL.scala 253:22]
  wire  s_2_322 = m_1747_io_s; // @[MUL.scala 252:21]
  wire  c_1_322 = m_1747_io_cout; // @[MUL.scala 253:22]
  wire  s_0_394 = m_1748_io_s; // @[MUL.scala 252:21]
  wire  c_0_394 = m_1748_io_cout; // @[MUL.scala 253:22]
  wire  s_2_323 = m_1749_io_s; // @[MUL.scala 252:21]
  wire  c_1_323 = m_1749_io_cout; // @[MUL.scala 253:22]
  wire  s_0_395 = m_1750_io_s; // @[MUL.scala 252:21]
  wire  c_0_395 = m_1750_io_cout; // @[MUL.scala 253:22]
  wire  s_2_324 = m_1751_io_s; // @[MUL.scala 252:21]
  wire  c_1_324 = m_1751_io_cout; // @[MUL.scala 253:22]
  wire  s_0_396 = m_1752_io_s; // @[MUL.scala 252:21]
  wire  c_0_396 = m_1752_io_cout; // @[MUL.scala 253:22]
  wire  s_2_325 = m_1753_io_s; // @[MUL.scala 252:21]
  wire  c_1_325 = m_1753_io_cout; // @[MUL.scala 253:22]
  wire  s_0_397 = m_1754_io_s; // @[MUL.scala 252:21]
  wire  c_0_397 = m_1754_io_cout; // @[MUL.scala 253:22]
  wire  s_2_326 = m_1755_io_s; // @[MUL.scala 252:21]
  wire  c_1_326 = m_1755_io_cout; // @[MUL.scala 253:22]
  wire  s_0_398 = m_1756_io_s; // @[MUL.scala 252:21]
  wire  c_0_398 = m_1756_io_cout; // @[MUL.scala 253:22]
  wire  s_2_327 = m_1757_io_s; // @[MUL.scala 252:21]
  wire  c_1_327 = m_1757_io_cout; // @[MUL.scala 253:22]
  wire  s_0_399 = m_1758_io_s; // @[MUL.scala 252:21]
  wire  c_0_399 = m_1758_io_cout; // @[MUL.scala 253:22]
  wire  s_2_328 = m_1759_io_s; // @[MUL.scala 252:21]
  wire  c_1_328 = m_1759_io_cout; // @[MUL.scala 253:22]
  wire  s_0_400 = m_1761_io_s; // @[MUL.scala 252:21]
  wire  c_0_400 = m_1761_io_cout; // @[MUL.scala 253:22]
  wire  s_2_329 = m_1762_io_s; // @[MUL.scala 252:21]
  wire  c_1_329 = m_1762_io_cout; // @[MUL.scala 253:22]
  wire  s_0_401 = m_1764_io_s; // @[MUL.scala 252:21]
  wire  c_0_401 = m_1764_io_cout; // @[MUL.scala 253:22]
  wire  s_2_330 = m_1765_io_s; // @[MUL.scala 252:21]
  wire  c_1_330 = m_1765_io_cout; // @[MUL.scala 253:22]
  wire  s_0_402 = m_1767_io_s; // @[MUL.scala 252:21]
  wire  c_0_402 = m_1767_io_cout; // @[MUL.scala 253:22]
  wire  s_2_331 = m_1768_io_s; // @[MUL.scala 252:21]
  wire  c_1_331 = m_1768_io_cout; // @[MUL.scala 253:22]
  wire  s_0_403 = m_1770_io_s; // @[MUL.scala 252:21]
  wire  c_0_403 = m_1770_io_cout; // @[MUL.scala 253:22]
  wire  s_2_332 = m_1771_io_s; // @[MUL.scala 252:21]
  wire  c_1_332 = m_1771_io_cout; // @[MUL.scala 253:22]
  wire  s_0_404 = m_1773_io_s; // @[MUL.scala 252:21]
  wire  c_0_404 = m_1773_io_cout; // @[MUL.scala 253:22]
  wire  s_2_333 = m_1774_io_s; // @[MUL.scala 252:21]
  wire  c_1_333 = m_1774_io_cout; // @[MUL.scala 253:22]
  wire  s_0_405 = m_1776_io_s; // @[MUL.scala 252:21]
  wire  c_0_405 = m_1776_io_cout; // @[MUL.scala 253:22]
  wire  s_2_334 = m_1777_io_s; // @[MUL.scala 252:21]
  wire  c_1_334 = m_1777_io_cout; // @[MUL.scala 253:22]
  wire  s_0_406 = m_1779_io_s; // @[MUL.scala 252:21]
  wire  c_0_406 = m_1779_io_cout; // @[MUL.scala 253:22]
  wire  s_2_335 = m_1780_io_s; // @[MUL.scala 252:21]
  wire  c_1_335 = m_1780_io_cout; // @[MUL.scala 253:22]
  wire  s_0_407 = m_1782_io_s; // @[MUL.scala 252:21]
  wire  c_0_407 = m_1782_io_cout; // @[MUL.scala 253:22]
  wire  s_2_336 = m_1783_io_s; // @[MUL.scala 252:21]
  wire  c_1_336 = m_1783_io_cout; // @[MUL.scala 253:22]
  wire  s_4_250 = m_1784_io_s; // @[MUL.scala 252:21]
  wire  c_2_250 = m_1784_io_cout; // @[MUL.scala 253:22]
  wire  s_0_408 = m_1785_io_s; // @[MUL.scala 252:21]
  wire  c_0_408 = m_1785_io_cout; // @[MUL.scala 253:22]
  wire  s_2_337 = m_1786_io_s; // @[MUL.scala 252:21]
  wire  c_1_337 = m_1786_io_cout; // @[MUL.scala 253:22]
  wire  s_4_251 = m_1787_io_s; // @[MUL.scala 252:21]
  wire  c_2_251 = m_1787_io_cout; // @[MUL.scala 253:22]
  wire  s_0_409 = m_1788_io_s; // @[MUL.scala 252:21]
  wire  c_0_409 = m_1788_io_cout; // @[MUL.scala 253:22]
  wire  s_2_338 = m_1789_io_s; // @[MUL.scala 252:21]
  wire  c_1_338 = m_1789_io_cout; // @[MUL.scala 253:22]
  wire  s_4_252 = m_1790_io_s; // @[MUL.scala 252:21]
  wire  c_2_252 = m_1790_io_cout; // @[MUL.scala 253:22]
  wire  s_0_410 = m_1791_io_s; // @[MUL.scala 252:21]
  wire  c_0_410 = m_1791_io_cout; // @[MUL.scala 253:22]
  wire  s_2_339 = m_1792_io_s; // @[MUL.scala 252:21]
  wire  c_1_339 = m_1792_io_cout; // @[MUL.scala 253:22]
  wire  s_4_253 = m_1793_io_s; // @[MUL.scala 252:21]
  wire  c_2_253 = m_1793_io_cout; // @[MUL.scala 253:22]
  wire  s_0_411 = m_1794_io_s; // @[MUL.scala 252:21]
  wire  c_0_411 = m_1794_io_cout; // @[MUL.scala 253:22]
  wire  s_2_340 = m_1795_io_s; // @[MUL.scala 252:21]
  wire  c_1_340 = m_1795_io_cout; // @[MUL.scala 253:22]
  wire  s_4_254 = m_1796_io_s; // @[MUL.scala 252:21]
  wire  c_2_254 = m_1796_io_cout; // @[MUL.scala 253:22]
  wire  s_0_412 = m_1797_io_s; // @[MUL.scala 252:21]
  wire  c_0_412 = m_1797_io_cout; // @[MUL.scala 253:22]
  wire  s_2_341 = m_1798_io_s; // @[MUL.scala 252:21]
  wire  c_1_341 = m_1798_io_cout; // @[MUL.scala 253:22]
  wire  s_4_255 = m_1799_io_s; // @[MUL.scala 252:21]
  wire  c_2_255 = m_1799_io_cout; // @[MUL.scala 253:22]
  wire  s_0_413 = m_1800_io_s; // @[MUL.scala 252:21]
  wire  c_0_413 = m_1800_io_cout; // @[MUL.scala 253:22]
  wire  s_2_342 = m_1801_io_s; // @[MUL.scala 252:21]
  wire  c_1_342 = m_1801_io_cout; // @[MUL.scala 253:22]
  wire  s_4_256 = m_1802_io_s; // @[MUL.scala 252:21]
  wire  c_2_256 = m_1802_io_cout; // @[MUL.scala 253:22]
  wire  s_0_414 = m_1803_io_s; // @[MUL.scala 252:21]
  wire  c_0_414 = m_1803_io_cout; // @[MUL.scala 253:22]
  wire  s_2_343 = m_1804_io_s; // @[MUL.scala 252:21]
  wire  c_1_343 = m_1804_io_cout; // @[MUL.scala 253:22]
  wire  s_4_257 = m_1805_io_s; // @[MUL.scala 252:21]
  wire  c_2_257 = m_1805_io_cout; // @[MUL.scala 253:22]
  wire  s_0_415 = m_1806_io_s; // @[MUL.scala 252:21]
  wire  c_0_415 = m_1806_io_cout; // @[MUL.scala 253:22]
  wire  s_2_344 = m_1807_io_s; // @[MUL.scala 252:21]
  wire  c_1_344 = m_1807_io_cout; // @[MUL.scala 253:22]
  wire  s_4_258 = m_1808_io_s; // @[MUL.scala 252:21]
  wire  c_2_258 = m_1808_io_cout; // @[MUL.scala 253:22]
  wire  s_0_416 = m_1809_io_s; // @[MUL.scala 252:21]
  wire  c_0_416 = m_1809_io_cout; // @[MUL.scala 253:22]
  wire  s_2_345 = m_1810_io_s; // @[MUL.scala 252:21]
  wire  c_1_345 = m_1810_io_cout; // @[MUL.scala 253:22]
  wire  s_4_259 = m_1811_io_s; // @[MUL.scala 252:21]
  wire  c_2_259 = m_1811_io_cout; // @[MUL.scala 253:22]
  wire  s_0_417 = m_1812_io_s; // @[MUL.scala 252:21]
  wire  c_0_417 = m_1812_io_cout; // @[MUL.scala 253:22]
  wire  s_2_346 = m_1813_io_s; // @[MUL.scala 252:21]
  wire  c_1_346 = m_1813_io_cout; // @[MUL.scala 253:22]
  wire  s_4_260 = m_1814_io_s; // @[MUL.scala 252:21]
  wire  c_2_260 = m_1814_io_cout; // @[MUL.scala 253:22]
  wire  s_0_418 = m_1815_io_s; // @[MUL.scala 252:21]
  wire  c_0_418 = m_1815_io_cout; // @[MUL.scala 253:22]
  wire  s_2_347 = m_1816_io_s; // @[MUL.scala 252:21]
  wire  c_1_347 = m_1816_io_cout; // @[MUL.scala 253:22]
  wire  s_4_261 = m_1817_io_s; // @[MUL.scala 252:21]
  wire  c_2_261 = m_1817_io_cout; // @[MUL.scala 253:22]
  wire  s_0_419 = m_1818_io_s; // @[MUL.scala 252:21]
  wire  c_0_419 = m_1818_io_cout; // @[MUL.scala 253:22]
  wire  s_2_348 = m_1819_io_s; // @[MUL.scala 252:21]
  wire  c_1_348 = m_1819_io_cout; // @[MUL.scala 253:22]
  wire  s_4_262 = m_1820_io_s; // @[MUL.scala 252:21]
  wire  c_2_262 = m_1820_io_cout; // @[MUL.scala 253:22]
  wire  s_0_420 = m_1821_io_s; // @[MUL.scala 252:21]
  wire  c_0_420 = m_1821_io_cout; // @[MUL.scala 253:22]
  wire  s_2_349 = m_1822_io_s; // @[MUL.scala 252:21]
  wire  c_1_349 = m_1822_io_cout; // @[MUL.scala 253:22]
  wire  s_4_263 = m_1823_io_s; // @[MUL.scala 252:21]
  wire  c_2_263 = m_1823_io_cout; // @[MUL.scala 253:22]
  wire  s_0_421 = m_1824_io_s; // @[MUL.scala 252:21]
  wire  c_0_421 = m_1824_io_cout; // @[MUL.scala 253:22]
  wire  s_2_350 = m_1825_io_s; // @[MUL.scala 252:21]
  wire  c_1_350 = m_1825_io_cout; // @[MUL.scala 253:22]
  wire  s_4_264 = m_1826_io_s; // @[MUL.scala 252:21]
  wire  c_2_264 = m_1826_io_cout; // @[MUL.scala 253:22]
  wire  s_0_422 = m_1827_io_s; // @[MUL.scala 252:21]
  wire  c_0_422 = m_1827_io_cout; // @[MUL.scala 253:22]
  wire  s_2_351 = m_1828_io_s; // @[MUL.scala 252:21]
  wire  c_1_351 = m_1828_io_cout; // @[MUL.scala 253:22]
  wire  s_4_265 = m_1829_io_s; // @[MUL.scala 252:21]
  wire  c_2_265 = m_1829_io_cout; // @[MUL.scala 253:22]
  wire  s_0_423 = m_1830_io_s; // @[MUL.scala 252:21]
  wire  c_0_423 = m_1830_io_cout; // @[MUL.scala 253:22]
  wire  s_2_352 = m_1831_io_s; // @[MUL.scala 252:21]
  wire  c_1_352 = m_1831_io_cout; // @[MUL.scala 253:22]
  wire  s_4_266 = m_1832_io_s; // @[MUL.scala 252:21]
  wire  c_2_266 = m_1832_io_cout; // @[MUL.scala 253:22]
  wire  s_0_424 = m_1833_io_s; // @[MUL.scala 252:21]
  wire  c_0_424 = m_1833_io_cout; // @[MUL.scala 253:22]
  wire  s_2_353 = m_1834_io_s; // @[MUL.scala 252:21]
  wire  c_1_353 = m_1834_io_cout; // @[MUL.scala 253:22]
  wire  s_4_267 = m_1835_io_s; // @[MUL.scala 252:21]
  wire  c_2_267 = m_1835_io_cout; // @[MUL.scala 253:22]
  wire  s_0_425 = m_1836_io_s; // @[MUL.scala 252:21]
  wire  c_0_425 = m_1836_io_cout; // @[MUL.scala 253:22]
  wire  s_2_354 = m_1837_io_s; // @[MUL.scala 252:21]
  wire  c_1_354 = m_1837_io_cout; // @[MUL.scala 253:22]
  wire  s_4_268 = m_1838_io_s; // @[MUL.scala 252:21]
  wire  c_2_268 = m_1838_io_cout; // @[MUL.scala 253:22]
  wire  s_0_426 = m_1839_io_s; // @[MUL.scala 252:21]
  wire  c_0_426 = m_1839_io_cout; // @[MUL.scala 253:22]
  wire  s_2_355 = m_1840_io_s; // @[MUL.scala 252:21]
  wire  c_1_355 = m_1840_io_cout; // @[MUL.scala 253:22]
  wire  s_4_269 = m_1841_io_s; // @[MUL.scala 252:21]
  wire  c_2_269 = m_1841_io_cout; // @[MUL.scala 253:22]
  wire  s_0_427 = m_1842_io_s; // @[MUL.scala 252:21]
  wire  c_0_427 = m_1842_io_cout; // @[MUL.scala 253:22]
  wire  s_2_356 = m_1843_io_s; // @[MUL.scala 252:21]
  wire  c_1_356 = m_1843_io_cout; // @[MUL.scala 253:22]
  wire  s_4_270 = m_1844_io_s; // @[MUL.scala 252:21]
  wire  c_2_270 = m_1844_io_cout; // @[MUL.scala 253:22]
  wire  s_0_428 = m_1845_io_s; // @[MUL.scala 252:21]
  wire  c_0_428 = m_1845_io_cout; // @[MUL.scala 253:22]
  wire  s_2_357 = m_1846_io_s; // @[MUL.scala 252:21]
  wire  c_1_357 = m_1846_io_cout; // @[MUL.scala 253:22]
  wire  s_4_271 = m_1847_io_s; // @[MUL.scala 252:21]
  wire  c_2_271 = m_1847_io_cout; // @[MUL.scala 253:22]
  wire  s_0_429 = m_1848_io_s; // @[MUL.scala 252:21]
  wire  c_0_429 = m_1848_io_cout; // @[MUL.scala 253:22]
  wire  s_2_358 = m_1849_io_s; // @[MUL.scala 252:21]
  wire  c_1_358 = m_1849_io_cout; // @[MUL.scala 253:22]
  wire  s_4_272 = m_1850_io_s; // @[MUL.scala 252:21]
  wire  c_2_272 = m_1850_io_cout; // @[MUL.scala 253:22]
  wire  s_0_430 = m_1851_io_s; // @[MUL.scala 252:21]
  wire  c_0_430 = m_1851_io_cout; // @[MUL.scala 253:22]
  wire  s_2_359 = m_1852_io_s; // @[MUL.scala 252:21]
  wire  c_1_359 = m_1852_io_cout; // @[MUL.scala 253:22]
  wire  s_4_273 = m_1853_io_s; // @[MUL.scala 252:21]
  wire  c_2_273 = m_1853_io_cout; // @[MUL.scala 253:22]
  wire  s_0_431 = m_1854_io_s; // @[MUL.scala 252:21]
  wire  c_0_431 = m_1854_io_cout; // @[MUL.scala 253:22]
  wire  s_2_360 = m_1855_io_s; // @[MUL.scala 252:21]
  wire  c_1_360 = m_1855_io_cout; // @[MUL.scala 253:22]
  wire  s_4_274 = m_1856_io_s; // @[MUL.scala 252:21]
  wire  c_2_274 = m_1856_io_cout; // @[MUL.scala 253:22]
  wire  s_0_432 = m_1857_io_s; // @[MUL.scala 252:21]
  wire  c_0_432 = m_1857_io_cout; // @[MUL.scala 253:22]
  wire  s_2_361 = m_1858_io_s; // @[MUL.scala 252:21]
  wire  c_1_361 = m_1858_io_cout; // @[MUL.scala 253:22]
  wire  s_4_275 = m_1859_io_s; // @[MUL.scala 252:21]
  wire  c_2_275 = m_1859_io_cout; // @[MUL.scala 253:22]
  wire  s_0_433 = m_1860_io_s; // @[MUL.scala 252:21]
  wire  c_0_433 = m_1860_io_cout; // @[MUL.scala 253:22]
  wire  s_2_362 = m_1861_io_s; // @[MUL.scala 252:21]
  wire  c_1_362 = m_1861_io_cout; // @[MUL.scala 253:22]
  wire  s_4_276 = m_1862_io_s; // @[MUL.scala 252:21]
  wire  c_2_276 = m_1862_io_cout; // @[MUL.scala 253:22]
  wire  s_0_434 = m_1863_io_s; // @[MUL.scala 252:21]
  wire  c_0_434 = m_1863_io_cout; // @[MUL.scala 253:22]
  wire  s_2_363 = m_1864_io_s; // @[MUL.scala 252:21]
  wire  c_1_363 = m_1864_io_cout; // @[MUL.scala 253:22]
  wire  s_0_435 = m_1866_io_s; // @[MUL.scala 252:21]
  wire  c_0_435 = m_1866_io_cout; // @[MUL.scala 253:22]
  wire  s_2_364 = m_1867_io_s; // @[MUL.scala 252:21]
  wire  c_1_364 = m_1867_io_cout; // @[MUL.scala 253:22]
  wire  s_0_436 = m_1869_io_s; // @[MUL.scala 252:21]
  wire  c_0_436 = m_1869_io_cout; // @[MUL.scala 253:22]
  wire  s_2_365 = m_1870_io_s; // @[MUL.scala 252:21]
  wire  c_1_365 = m_1870_io_cout; // @[MUL.scala 253:22]
  wire  s_0_437 = m_1872_io_s; // @[MUL.scala 252:21]
  wire  c_0_437 = m_1872_io_cout; // @[MUL.scala 253:22]
  wire  s_2_366 = m_1873_io_s; // @[MUL.scala 252:21]
  wire  c_1_366 = m_1873_io_cout; // @[MUL.scala 253:22]
  wire  s_0_438 = m_1875_io_s; // @[MUL.scala 252:21]
  wire  c_0_438 = m_1875_io_cout; // @[MUL.scala 253:22]
  wire  s_2_367 = m_1876_io_s; // @[MUL.scala 252:21]
  wire  c_1_367 = m_1876_io_cout; // @[MUL.scala 253:22]
  wire  s_0_439 = m_1878_io_s; // @[MUL.scala 252:21]
  wire  c_0_439 = m_1878_io_cout; // @[MUL.scala 253:22]
  wire  s_2_368 = m_1879_io_s; // @[MUL.scala 252:21]
  wire  c_1_368 = m_1879_io_cout; // @[MUL.scala 253:22]
  wire  s_0_440 = m_1881_io_s; // @[MUL.scala 252:21]
  wire  c_0_440 = m_1881_io_cout; // @[MUL.scala 253:22]
  wire  s_2_369 = m_1882_io_s; // @[MUL.scala 252:21]
  wire  c_1_369 = m_1882_io_cout; // @[MUL.scala 253:22]
  wire  s_0_441 = m_1884_io_s; // @[MUL.scala 252:21]
  wire  c_0_441 = m_1884_io_cout; // @[MUL.scala 253:22]
  wire  s_2_370 = m_1885_io_s; // @[MUL.scala 252:21]
  wire  c_1_370 = m_1885_io_cout; // @[MUL.scala 253:22]
  wire  s_0_442 = m_1887_io_s; // @[MUL.scala 252:21]
  wire  c_0_442 = m_1887_io_cout; // @[MUL.scala 253:22]
  wire  s_2_371 = m_1888_io_s; // @[MUL.scala 252:21]
  wire  c_1_371 = m_1888_io_cout; // @[MUL.scala 253:22]
  wire  s_0_443 = m_1890_io_s; // @[MUL.scala 252:21]
  wire  c_0_443 = m_1890_io_cout; // @[MUL.scala 253:22]
  wire  s_2_372 = m_1891_io_s; // @[MUL.scala 252:21]
  wire  c_1_372 = m_1891_io_cout; // @[MUL.scala 253:22]
  wire  s_0_444 = m_1893_io_s; // @[MUL.scala 252:21]
  wire  c_0_444 = m_1893_io_cout; // @[MUL.scala 253:22]
  wire  s_2_373 = m_1894_io_s; // @[MUL.scala 252:21]
  wire  c_1_373 = m_1894_io_cout; // @[MUL.scala 253:22]
  wire  s_0_445 = m_1896_io_s; // @[MUL.scala 252:21]
  wire  c_0_445 = m_1896_io_cout; // @[MUL.scala 253:22]
  wire  s_2_374 = m_1897_io_s; // @[MUL.scala 252:21]
  wire  c_1_374 = m_1897_io_cout; // @[MUL.scala 253:22]
  wire  s_0_446 = m_1898_io_s; // @[MUL.scala 252:21]
  wire  c_0_446 = m_1898_io_cout; // @[MUL.scala 253:22]
  wire  s_2_375 = m_1899_io_s; // @[MUL.scala 252:21]
  wire  c_1_375 = m_1899_io_cout; // @[MUL.scala 253:22]
  wire  s_0_447 = m_1900_io_s; // @[MUL.scala 252:21]
  wire  c_0_447 = m_1900_io_cout; // @[MUL.scala 253:22]
  wire  s_2_376 = m_1901_io_s; // @[MUL.scala 252:21]
  wire  c_1_376 = m_1901_io_cout; // @[MUL.scala 253:22]
  wire  s_0_448 = m_1902_io_s; // @[MUL.scala 252:21]
  wire  c_0_448 = m_1902_io_cout; // @[MUL.scala 253:22]
  wire  s_2_377 = m_1903_io_s; // @[MUL.scala 252:21]
  wire  c_1_377 = m_1903_io_cout; // @[MUL.scala 253:22]
  wire  s_0_449 = m_1904_io_s; // @[MUL.scala 252:21]
  wire  c_0_449 = m_1904_io_cout; // @[MUL.scala 253:22]
  wire  s_2_378 = m_1905_io_s; // @[MUL.scala 252:21]
  wire  c_1_378 = m_1905_io_cout; // @[MUL.scala 253:22]
  wire  s_0_450 = m_1906_io_s; // @[MUL.scala 252:21]
  wire  c_0_450 = m_1906_io_cout; // @[MUL.scala 253:22]
  wire  s_2_379 = m_1907_io_s; // @[MUL.scala 252:21]
  wire  c_1_379 = m_1907_io_cout; // @[MUL.scala 253:22]
  wire  s_0_451 = m_1908_io_s; // @[MUL.scala 252:21]
  wire  c_0_451 = m_1908_io_cout; // @[MUL.scala 253:22]
  wire  s_2_380 = m_1909_io_s; // @[MUL.scala 252:21]
  wire  c_1_380 = m_1909_io_cout; // @[MUL.scala 253:22]
  wire  s_0_452 = m_1910_io_s; // @[MUL.scala 252:21]
  wire  c_0_452 = m_1910_io_cout; // @[MUL.scala 253:22]
  wire  s_2_381 = m_1911_io_s; // @[MUL.scala 252:21]
  wire  c_1_381 = m_1911_io_cout; // @[MUL.scala 253:22]
  wire  s_0_453 = m_1912_io_s; // @[MUL.scala 252:21]
  wire  c_0_453 = m_1912_io_cout; // @[MUL.scala 253:22]
  wire  s_2_382 = m_1913_io_s; // @[MUL.scala 252:21]
  wire  c_1_382 = m_1913_io_cout; // @[MUL.scala 253:22]
  wire  s_0_454 = m_1914_io_s; // @[MUL.scala 252:21]
  wire  c_0_454 = m_1914_io_cout; // @[MUL.scala 253:22]
  wire  s_2_383 = m_1915_io_s; // @[MUL.scala 252:21]
  wire  c_1_383 = m_1915_io_cout; // @[MUL.scala 253:22]
  wire  s_0_455 = m_1916_io_s; // @[MUL.scala 252:21]
  wire  c_0_455 = m_1916_io_cout; // @[MUL.scala 253:22]
  wire  s_2_384 = m_1917_io_s; // @[MUL.scala 252:21]
  wire  c_1_384 = m_1917_io_cout; // @[MUL.scala 253:22]
  wire  s_0_456 = m_1918_io_s; // @[MUL.scala 252:21]
  wire  c_0_456 = m_1918_io_cout; // @[MUL.scala 253:22]
  wire  s_2_385 = m_1919_io_s; // @[MUL.scala 252:21]
  wire  c_1_385 = m_1919_io_cout; // @[MUL.scala 253:22]
  wire  s_0_457 = m_1920_io_s; // @[MUL.scala 252:21]
  wire  c_0_457 = m_1920_io_cout; // @[MUL.scala 253:22]
  wire  s_2_386 = m_1921_io_s; // @[MUL.scala 252:21]
  wire  c_1_386 = m_1921_io_cout; // @[MUL.scala 253:22]
  wire  s_0_458 = m_1922_io_s; // @[MUL.scala 252:21]
  wire  c_0_458 = m_1922_io_cout; // @[MUL.scala 253:22]
  wire  s_2_387 = m_1923_io_s; // @[MUL.scala 252:21]
  wire  c_1_387 = m_1923_io_cout; // @[MUL.scala 253:22]
  wire  s_0_459 = m_1924_io_s; // @[MUL.scala 252:21]
  wire  c_0_459 = m_1924_io_cout; // @[MUL.scala 253:22]
  wire  s_0_460 = m_1926_io_s; // @[MUL.scala 252:21]
  wire  c_0_460 = m_1926_io_cout; // @[MUL.scala 253:22]
  wire  s_0_461 = m_1928_io_s; // @[MUL.scala 252:21]
  wire  c_0_461 = m_1928_io_cout; // @[MUL.scala 253:22]
  wire  s_0_462 = m_1930_io_s; // @[MUL.scala 252:21]
  wire  c_0_462 = m_1930_io_cout; // @[MUL.scala 253:22]
  wire  s_0_463 = m_1931_io_s; // @[MUL.scala 252:21]
  wire  c_0_463 = m_1931_io_cout; // @[MUL.scala 253:22]
  wire  s_0_464 = m_1932_io_s; // @[MUL.scala 252:21]
  wire  c_0_464 = m_1932_io_cout; // @[MUL.scala 253:22]
  wire  s_0_465 = m_1933_io_s; // @[MUL.scala 252:21]
  wire  c_0_465 = m_1933_io_cout; // @[MUL.scala 253:22]
  wire  s_0_466 = m_1934_io_s; // @[MUL.scala 252:21]
  wire  c_0_466 = m_1934_io_cout; // @[MUL.scala 253:22]
  wire  s_0_467 = m_1935_io_s; // @[MUL.scala 252:21]
  wire  c_0_467 = m_1935_io_cout; // @[MUL.scala 253:22]
  wire  s_0_468 = m_1936_io_s; // @[MUL.scala 252:21]
  wire  c_0_468 = m_1936_io_cout; // @[MUL.scala 253:22]
  wire  s_0_469 = m_1937_io_s; // @[MUL.scala 252:21]
  wire  c_0_469 = m_1937_io_cout; // @[MUL.scala 253:22]
  wire  s_0_470 = m_1938_io_s; // @[MUL.scala 252:21]
  wire  c_0_470 = m_1938_io_cout; // @[MUL.scala 253:22]
  wire  s_0_471 = m_1939_io_s; // @[MUL.scala 252:21]
  wire  c_0_471 = m_1939_io_cout; // @[MUL.scala 253:22]
  wire  s_0_472 = m_1940_io_s; // @[MUL.scala 252:21]
  wire  c_0_472 = m_1940_io_cout; // @[MUL.scala 253:22]
  wire  s_0_473 = m_1941_io_s; // @[MUL.scala 252:21]
  wire  c_0_473 = m_1941_io_cout; // @[MUL.scala 253:22]
  wire  s_0_474 = m_1942_io_s; // @[MUL.scala 252:21]
  wire  c_0_474 = m_1942_io_cout; // @[MUL.scala 253:22]
  wire  s_0_475 = m_1943_io_s; // @[MUL.scala 252:21]
  wire  c_0_475 = m_1943_io_cout; // @[MUL.scala 253:22]
  reg  r_2308; // @[Reg.scala 16:16]
  reg  r_2309; // @[Reg.scala 16:16]
  reg  r_2310; // @[Reg.scala 16:16]
  reg  r_2311; // @[Reg.scala 16:16]
  reg  r_2312; // @[Reg.scala 16:16]
  reg  r_2313; // @[Reg.scala 16:16]
  reg  r_2314; // @[Reg.scala 16:16]
  reg  r_2315; // @[Reg.scala 16:16]
  reg  r_2316; // @[Reg.scala 16:16]
  reg  r_2317; // @[Reg.scala 16:16]
  reg  r_2318; // @[Reg.scala 16:16]
  reg  r_2319; // @[Reg.scala 16:16]
  reg  r_2320; // @[Reg.scala 16:16]
  reg  r_2321; // @[Reg.scala 16:16]
  reg  r_2322; // @[Reg.scala 16:16]
  reg  r_2323; // @[Reg.scala 16:16]
  reg  r_2324; // @[Reg.scala 16:16]
  reg  r_2325; // @[Reg.scala 16:16]
  reg  r_2326; // @[Reg.scala 16:16]
  reg  r_2327; // @[Reg.scala 16:16]
  reg  r_2328; // @[Reg.scala 16:16]
  reg  r_2329; // @[Reg.scala 16:16]
  reg  r_2330; // @[Reg.scala 16:16]
  reg  r_2331; // @[Reg.scala 16:16]
  reg  r_2332; // @[Reg.scala 16:16]
  reg  r_2333; // @[Reg.scala 16:16]
  reg  r_2334; // @[Reg.scala 16:16]
  reg  r_2335; // @[Reg.scala 16:16]
  reg  r_2336; // @[Reg.scala 16:16]
  reg  r_2337; // @[Reg.scala 16:16]
  reg  r_2338; // @[Reg.scala 16:16]
  reg  r_2339; // @[Reg.scala 16:16]
  reg  r_2340; // @[Reg.scala 16:16]
  reg  r_2341; // @[Reg.scala 16:16]
  reg  r_2342; // @[Reg.scala 16:16]
  reg  r_2343; // @[Reg.scala 16:16]
  reg  r_2344; // @[Reg.scala 16:16]
  reg  r_2345; // @[Reg.scala 16:16]
  reg  r_2346; // @[Reg.scala 16:16]
  reg  r_2347; // @[Reg.scala 16:16]
  reg  r_2348; // @[Reg.scala 16:16]
  reg  r_2349; // @[Reg.scala 16:16]
  reg  r_2350; // @[Reg.scala 16:16]
  reg  r_2351; // @[Reg.scala 16:16]
  reg  r_2352; // @[Reg.scala 16:16]
  reg  r_2353; // @[Reg.scala 16:16]
  reg  r_2354; // @[Reg.scala 16:16]
  reg  r_2355; // @[Reg.scala 16:16]
  reg  r_2356; // @[Reg.scala 16:16]
  reg  r_2357; // @[Reg.scala 16:16]
  reg  r_2358; // @[Reg.scala 16:16]
  reg  r_2359; // @[Reg.scala 16:16]
  reg  r_2360; // @[Reg.scala 16:16]
  reg  r_2361; // @[Reg.scala 16:16]
  reg  r_2362; // @[Reg.scala 16:16]
  reg  r_2363; // @[Reg.scala 16:16]
  reg  r_2364; // @[Reg.scala 16:16]
  reg  r_2365; // @[Reg.scala 16:16]
  reg  r_2366; // @[Reg.scala 16:16]
  reg  r_2367; // @[Reg.scala 16:16]
  reg  r_2368; // @[Reg.scala 16:16]
  reg  r_2369; // @[Reg.scala 16:16]
  reg  r_2370; // @[Reg.scala 16:16]
  reg  r_2371; // @[Reg.scala 16:16]
  reg  r_2372; // @[Reg.scala 16:16]
  reg  r_2373; // @[Reg.scala 16:16]
  reg  r_2374; // @[Reg.scala 16:16]
  reg  r_2375; // @[Reg.scala 16:16]
  reg  r_2376; // @[Reg.scala 16:16]
  reg  r_2377; // @[Reg.scala 16:16]
  reg  r_2378; // @[Reg.scala 16:16]
  reg  r_2379; // @[Reg.scala 16:16]
  reg  r_2380; // @[Reg.scala 16:16]
  reg  r_2381; // @[Reg.scala 16:16]
  reg  r_2382; // @[Reg.scala 16:16]
  reg  r_2383; // @[Reg.scala 16:16]
  reg  r_2384; // @[Reg.scala 16:16]
  reg  r_2385; // @[Reg.scala 16:16]
  reg  r_2386; // @[Reg.scala 16:16]
  reg  r_2387; // @[Reg.scala 16:16]
  reg  r_2388; // @[Reg.scala 16:16]
  reg  r_2389; // @[Reg.scala 16:16]
  reg  r_2390; // @[Reg.scala 16:16]
  reg  r_2391; // @[Reg.scala 16:16]
  reg  r_2392; // @[Reg.scala 16:16]
  reg  r_2393; // @[Reg.scala 16:16]
  reg  r_2394; // @[Reg.scala 16:16]
  reg  r_2395; // @[Reg.scala 16:16]
  reg  r_2396; // @[Reg.scala 16:16]
  reg  r_2397; // @[Reg.scala 16:16]
  reg  r_2398; // @[Reg.scala 16:16]
  reg  r_2399; // @[Reg.scala 16:16]
  reg  r_2400; // @[Reg.scala 16:16]
  reg  r_2401; // @[Reg.scala 16:16]
  reg  r_2402; // @[Reg.scala 16:16]
  reg  r_2403; // @[Reg.scala 16:16]
  reg  r_2404; // @[Reg.scala 16:16]
  reg  r_2405; // @[Reg.scala 16:16]
  reg  r_2406; // @[Reg.scala 16:16]
  reg  r_2407; // @[Reg.scala 16:16]
  reg  r_2408; // @[Reg.scala 16:16]
  reg  r_2409; // @[Reg.scala 16:16]
  reg  r_2410; // @[Reg.scala 16:16]
  reg  r_2411; // @[Reg.scala 16:16]
  reg  r_2412; // @[Reg.scala 16:16]
  reg  r_2413; // @[Reg.scala 16:16]
  reg  r_2414; // @[Reg.scala 16:16]
  reg  r_2415; // @[Reg.scala 16:16]
  reg  r_2416; // @[Reg.scala 16:16]
  reg  r_2417; // @[Reg.scala 16:16]
  reg  r_2418; // @[Reg.scala 16:16]
  reg  r_2419; // @[Reg.scala 16:16]
  reg  r_2420; // @[Reg.scala 16:16]
  reg  r_2421; // @[Reg.scala 16:16]
  reg  r_2422; // @[Reg.scala 16:16]
  reg  r_2423; // @[Reg.scala 16:16]
  reg  r_2424; // @[Reg.scala 16:16]
  reg  r_2425; // @[Reg.scala 16:16]
  reg  r_2426; // @[Reg.scala 16:16]
  reg  r_2427; // @[Reg.scala 16:16]
  reg  r_2428; // @[Reg.scala 16:16]
  reg  r_2429; // @[Reg.scala 16:16]
  reg  r_2430; // @[Reg.scala 16:16]
  reg  r_2431; // @[Reg.scala 16:16]
  reg  r_2432; // @[Reg.scala 16:16]
  reg  r_2433; // @[Reg.scala 16:16]
  reg  r_2434; // @[Reg.scala 16:16]
  reg  r_2435; // @[Reg.scala 16:16]
  reg  r_2436; // @[Reg.scala 16:16]
  reg  r_2437; // @[Reg.scala 16:16]
  reg  r_2438; // @[Reg.scala 16:16]
  reg  r_2439; // @[Reg.scala 16:16]
  reg  r_2440; // @[Reg.scala 16:16]
  reg  r_2441; // @[Reg.scala 16:16]
  reg  r_2442; // @[Reg.scala 16:16]
  reg  r_2443; // @[Reg.scala 16:16]
  reg  r_2444; // @[Reg.scala 16:16]
  reg  r_2445; // @[Reg.scala 16:16]
  reg  r_2446; // @[Reg.scala 16:16]
  reg  r_2447; // @[Reg.scala 16:16]
  reg  r_2448; // @[Reg.scala 16:16]
  reg  r_2449; // @[Reg.scala 16:16]
  reg  r_2450; // @[Reg.scala 16:16]
  reg  r_2451; // @[Reg.scala 16:16]
  reg  r_2452; // @[Reg.scala 16:16]
  reg  r_2453; // @[Reg.scala 16:16]
  reg  r_2454; // @[Reg.scala 16:16]
  reg  r_2455; // @[Reg.scala 16:16]
  reg  r_2456; // @[Reg.scala 16:16]
  reg  r_2457; // @[Reg.scala 16:16]
  reg  r_2458; // @[Reg.scala 16:16]
  reg  r_2459; // @[Reg.scala 16:16]
  reg  r_2460; // @[Reg.scala 16:16]
  reg  r_2461; // @[Reg.scala 16:16]
  reg  r_2462; // @[Reg.scala 16:16]
  reg  r_2463; // @[Reg.scala 16:16]
  reg  r_2464; // @[Reg.scala 16:16]
  reg  r_2465; // @[Reg.scala 16:16]
  reg  r_2466; // @[Reg.scala 16:16]
  reg  r_2467; // @[Reg.scala 16:16]
  reg  r_2468; // @[Reg.scala 16:16]
  reg  r_2469; // @[Reg.scala 16:16]
  reg  r_2470; // @[Reg.scala 16:16]
  reg  r_2471; // @[Reg.scala 16:16]
  reg  r_2472; // @[Reg.scala 16:16]
  reg  r_2473; // @[Reg.scala 16:16]
  reg  r_2474; // @[Reg.scala 16:16]
  reg  r_2475; // @[Reg.scala 16:16]
  reg  r_2476; // @[Reg.scala 16:16]
  reg  r_2477; // @[Reg.scala 16:16]
  reg  r_2478; // @[Reg.scala 16:16]
  reg  r_2479; // @[Reg.scala 16:16]
  reg  r_2480; // @[Reg.scala 16:16]
  reg  r_2481; // @[Reg.scala 16:16]
  reg  r_2482; // @[Reg.scala 16:16]
  reg  r_2483; // @[Reg.scala 16:16]
  reg  r_2484; // @[Reg.scala 16:16]
  reg  r_2485; // @[Reg.scala 16:16]
  reg  r_2486; // @[Reg.scala 16:16]
  reg  r_2487; // @[Reg.scala 16:16]
  reg  r_2488; // @[Reg.scala 16:16]
  reg  r_2489; // @[Reg.scala 16:16]
  reg  r_2490; // @[Reg.scala 16:16]
  reg  r_2491; // @[Reg.scala 16:16]
  reg  r_2492; // @[Reg.scala 16:16]
  reg  r_2493; // @[Reg.scala 16:16]
  reg  r_2494; // @[Reg.scala 16:16]
  reg  r_2495; // @[Reg.scala 16:16]
  reg  r_2496; // @[Reg.scala 16:16]
  reg  r_2497; // @[Reg.scala 16:16]
  reg  r_2498; // @[Reg.scala 16:16]
  reg  r_2499; // @[Reg.scala 16:16]
  reg  r_2500; // @[Reg.scala 16:16]
  reg  r_2501; // @[Reg.scala 16:16]
  reg  r_2502; // @[Reg.scala 16:16]
  reg  r_2503; // @[Reg.scala 16:16]
  reg  r_2504; // @[Reg.scala 16:16]
  reg  r_2505; // @[Reg.scala 16:16]
  reg  r_2506; // @[Reg.scala 16:16]
  reg  r_2507; // @[Reg.scala 16:16]
  reg  r_2508; // @[Reg.scala 16:16]
  reg  r_2509; // @[Reg.scala 16:16]
  reg  r_2510; // @[Reg.scala 16:16]
  reg  r_2511; // @[Reg.scala 16:16]
  reg  r_2512; // @[Reg.scala 16:16]
  reg  r_2513; // @[Reg.scala 16:16]
  reg  r_2514; // @[Reg.scala 16:16]
  reg  r_2515; // @[Reg.scala 16:16]
  reg  r_2516; // @[Reg.scala 16:16]
  reg  r_2517; // @[Reg.scala 16:16]
  reg  r_2518; // @[Reg.scala 16:16]
  reg  r_2519; // @[Reg.scala 16:16]
  reg  r_2520; // @[Reg.scala 16:16]
  reg  r_2521; // @[Reg.scala 16:16]
  reg  r_2522; // @[Reg.scala 16:16]
  reg  r_2523; // @[Reg.scala 16:16]
  reg  r_2524; // @[Reg.scala 16:16]
  reg  r_2525; // @[Reg.scala 16:16]
  reg  r_2526; // @[Reg.scala 16:16]
  reg  r_2527; // @[Reg.scala 16:16]
  reg  r_2528; // @[Reg.scala 16:16]
  reg  r_2529; // @[Reg.scala 16:16]
  reg  r_2530; // @[Reg.scala 16:16]
  reg  r_2531; // @[Reg.scala 16:16]
  reg  r_2532; // @[Reg.scala 16:16]
  reg  r_2533; // @[Reg.scala 16:16]
  reg  r_2534; // @[Reg.scala 16:16]
  reg  r_2535; // @[Reg.scala 16:16]
  reg  r_2536; // @[Reg.scala 16:16]
  reg  r_2537; // @[Reg.scala 16:16]
  reg  r_2538; // @[Reg.scala 16:16]
  reg  r_2539; // @[Reg.scala 16:16]
  reg  r_2540; // @[Reg.scala 16:16]
  reg  r_2541; // @[Reg.scala 16:16]
  reg  r_2542; // @[Reg.scala 16:16]
  reg  r_2543; // @[Reg.scala 16:16]
  reg  r_2544; // @[Reg.scala 16:16]
  reg  r_2545; // @[Reg.scala 16:16]
  reg  r_2546; // @[Reg.scala 16:16]
  reg  r_2547; // @[Reg.scala 16:16]
  reg  r_2548; // @[Reg.scala 16:16]
  reg  r_2549; // @[Reg.scala 16:16]
  reg  r_2550; // @[Reg.scala 16:16]
  reg  r_2551; // @[Reg.scala 16:16]
  reg  r_2552; // @[Reg.scala 16:16]
  reg  r_2553; // @[Reg.scala 16:16]
  reg  r_2554; // @[Reg.scala 16:16]
  reg  r_2555; // @[Reg.scala 16:16]
  reg  r_2556; // @[Reg.scala 16:16]
  reg  r_2557; // @[Reg.scala 16:16]
  reg  r_2558; // @[Reg.scala 16:16]
  reg  r_2559; // @[Reg.scala 16:16]
  reg  r_2560; // @[Reg.scala 16:16]
  reg  r_2561; // @[Reg.scala 16:16]
  reg  r_2562; // @[Reg.scala 16:16]
  reg  r_2563; // @[Reg.scala 16:16]
  reg  r_2564; // @[Reg.scala 16:16]
  reg  r_2565; // @[Reg.scala 16:16]
  reg  r_2566; // @[Reg.scala 16:16]
  reg  r_2567; // @[Reg.scala 16:16]
  reg  r_2568; // @[Reg.scala 16:16]
  reg  r_2569; // @[Reg.scala 16:16]
  reg  r_2570; // @[Reg.scala 16:16]
  reg  r_2571; // @[Reg.scala 16:16]
  reg  r_2572; // @[Reg.scala 16:16]
  reg  r_2573; // @[Reg.scala 16:16]
  reg  r_2574; // @[Reg.scala 16:16]
  reg  r_2575; // @[Reg.scala 16:16]
  reg  r_2576; // @[Reg.scala 16:16]
  reg  r_2577; // @[Reg.scala 16:16]
  reg  r_2578; // @[Reg.scala 16:16]
  reg  r_2579; // @[Reg.scala 16:16]
  reg  r_2580; // @[Reg.scala 16:16]
  reg  r_2581; // @[Reg.scala 16:16]
  reg  r_2582; // @[Reg.scala 16:16]
  reg  r_2583; // @[Reg.scala 16:16]
  reg  r_2584; // @[Reg.scala 16:16]
  reg  r_2585; // @[Reg.scala 16:16]
  reg  r_2586; // @[Reg.scala 16:16]
  reg  r_2587; // @[Reg.scala 16:16]
  reg  r_2588; // @[Reg.scala 16:16]
  reg  r_2589; // @[Reg.scala 16:16]
  reg  r_2590; // @[Reg.scala 16:16]
  reg  r_2591; // @[Reg.scala 16:16]
  reg  r_2592; // @[Reg.scala 16:16]
  reg  r_2593; // @[Reg.scala 16:16]
  reg  r_2594; // @[Reg.scala 16:16]
  reg  r_2595; // @[Reg.scala 16:16]
  reg  r_2596; // @[Reg.scala 16:16]
  reg  r_2597; // @[Reg.scala 16:16]
  reg  r_2598; // @[Reg.scala 16:16]
  reg  r_2599; // @[Reg.scala 16:16]
  reg  r_2600; // @[Reg.scala 16:16]
  reg  r_2601; // @[Reg.scala 16:16]
  reg  r_2602; // @[Reg.scala 16:16]
  reg  r_2603; // @[Reg.scala 16:16]
  reg  r_2604; // @[Reg.scala 16:16]
  reg  r_2605; // @[Reg.scala 16:16]
  reg  r_2606; // @[Reg.scala 16:16]
  reg  r_2607; // @[Reg.scala 16:16]
  reg  r_2608; // @[Reg.scala 16:16]
  reg  r_2609; // @[Reg.scala 16:16]
  reg  r_2610; // @[Reg.scala 16:16]
  reg  r_2611; // @[Reg.scala 16:16]
  reg  r_2612; // @[Reg.scala 16:16]
  reg  r_2613; // @[Reg.scala 16:16]
  reg  r_2614; // @[Reg.scala 16:16]
  reg  r_2615; // @[Reg.scala 16:16]
  reg  r_2616; // @[Reg.scala 16:16]
  reg  r_2617; // @[Reg.scala 16:16]
  reg  r_2618; // @[Reg.scala 16:16]
  reg  r_2619; // @[Reg.scala 16:16]
  reg  r_2620; // @[Reg.scala 16:16]
  reg  r_2621; // @[Reg.scala 16:16]
  reg  r_2622; // @[Reg.scala 16:16]
  reg  r_2623; // @[Reg.scala 16:16]
  reg  r_2624; // @[Reg.scala 16:16]
  reg  r_2625; // @[Reg.scala 16:16]
  reg  r_2626; // @[Reg.scala 16:16]
  reg  r_2627; // @[Reg.scala 16:16]
  reg  r_2628; // @[Reg.scala 16:16]
  reg  r_2629; // @[Reg.scala 16:16]
  reg  r_2630; // @[Reg.scala 16:16]
  reg  r_2631; // @[Reg.scala 16:16]
  reg  r_2632; // @[Reg.scala 16:16]
  reg  r_2633; // @[Reg.scala 16:16]
  reg  r_2634; // @[Reg.scala 16:16]
  reg  r_2635; // @[Reg.scala 16:16]
  reg  r_2636; // @[Reg.scala 16:16]
  reg  r_2637; // @[Reg.scala 16:16]
  reg  r_2638; // @[Reg.scala 16:16]
  reg  r_2639; // @[Reg.scala 16:16]
  reg  r_2640; // @[Reg.scala 16:16]
  reg  r_2641; // @[Reg.scala 16:16]
  reg  r_2642; // @[Reg.scala 16:16]
  reg  r_2643; // @[Reg.scala 16:16]
  reg  r_2644; // @[Reg.scala 16:16]
  reg  r_2645; // @[Reg.scala 16:16]
  reg  r_2646; // @[Reg.scala 16:16]
  reg  r_2647; // @[Reg.scala 16:16]
  reg  r_2648; // @[Reg.scala 16:16]
  reg  r_2649; // @[Reg.scala 16:16]
  reg  r_2650; // @[Reg.scala 16:16]
  reg  r_2651; // @[Reg.scala 16:16]
  reg  r_2652; // @[Reg.scala 16:16]
  reg  r_2653; // @[Reg.scala 16:16]
  reg  r_2654; // @[Reg.scala 16:16]
  reg  r_2655; // @[Reg.scala 16:16]
  reg  r_2656; // @[Reg.scala 16:16]
  reg  r_2657; // @[Reg.scala 16:16]
  reg  r_2658; // @[Reg.scala 16:16]
  reg  r_2659; // @[Reg.scala 16:16]
  reg  r_2660; // @[Reg.scala 16:16]
  reg  r_2661; // @[Reg.scala 16:16]
  reg  r_2662; // @[Reg.scala 16:16]
  reg  r_2663; // @[Reg.scala 16:16]
  reg  r_2664; // @[Reg.scala 16:16]
  reg  r_2665; // @[Reg.scala 16:16]
  reg  r_2666; // @[Reg.scala 16:16]
  reg  r_2667; // @[Reg.scala 16:16]
  reg  r_2668; // @[Reg.scala 16:16]
  reg  r_2669; // @[Reg.scala 16:16]
  reg  r_2670; // @[Reg.scala 16:16]
  reg  r_2671; // @[Reg.scala 16:16]
  reg  r_2672; // @[Reg.scala 16:16]
  reg  r_2673; // @[Reg.scala 16:16]
  reg  r_2674; // @[Reg.scala 16:16]
  reg  r_2675; // @[Reg.scala 16:16]
  reg  r_2676; // @[Reg.scala 16:16]
  reg  r_2677; // @[Reg.scala 16:16]
  reg  r_2678; // @[Reg.scala 16:16]
  reg  r_2679; // @[Reg.scala 16:16]
  reg  r_2680; // @[Reg.scala 16:16]
  reg  r_2681; // @[Reg.scala 16:16]
  reg  r_2682; // @[Reg.scala 16:16]
  reg  r_2683; // @[Reg.scala 16:16]
  reg  r_2684; // @[Reg.scala 16:16]
  reg  r_2685; // @[Reg.scala 16:16]
  reg  r_2686; // @[Reg.scala 16:16]
  reg  r_2687; // @[Reg.scala 16:16]
  reg  r_2688; // @[Reg.scala 16:16]
  reg  r_2689; // @[Reg.scala 16:16]
  reg  r_2690; // @[Reg.scala 16:16]
  reg  r_2691; // @[Reg.scala 16:16]
  reg  r_2692; // @[Reg.scala 16:16]
  reg  r_2693; // @[Reg.scala 16:16]
  reg  r_2694; // @[Reg.scala 16:16]
  reg  r_2695; // @[Reg.scala 16:16]
  reg  r_2696; // @[Reg.scala 16:16]
  reg  r_2697; // @[Reg.scala 16:16]
  reg  r_2698; // @[Reg.scala 16:16]
  reg  r_2699; // @[Reg.scala 16:16]
  reg  r_2700; // @[Reg.scala 16:16]
  reg  r_2701; // @[Reg.scala 16:16]
  reg  r_2702; // @[Reg.scala 16:16]
  reg  r_2703; // @[Reg.scala 16:16]
  reg  r_2704; // @[Reg.scala 16:16]
  reg  r_2705; // @[Reg.scala 16:16]
  reg  r_2706; // @[Reg.scala 16:16]
  reg  r_2707; // @[Reg.scala 16:16]
  reg  r_2708; // @[Reg.scala 16:16]
  reg  r_2709; // @[Reg.scala 16:16]
  reg  r_2710; // @[Reg.scala 16:16]
  reg  r_2711; // @[Reg.scala 16:16]
  reg  r_2712; // @[Reg.scala 16:16]
  reg  r_2713; // @[Reg.scala 16:16]
  reg  r_2714; // @[Reg.scala 16:16]
  reg  r_2715; // @[Reg.scala 16:16]
  reg  r_2716; // @[Reg.scala 16:16]
  reg  r_2717; // @[Reg.scala 16:16]
  reg  r_2718; // @[Reg.scala 16:16]
  reg  r_2719; // @[Reg.scala 16:16]
  reg  r_2720; // @[Reg.scala 16:16]
  reg  r_2721; // @[Reg.scala 16:16]
  reg  r_2722; // @[Reg.scala 16:16]
  reg  r_2723; // @[Reg.scala 16:16]
  reg  r_2724; // @[Reg.scala 16:16]
  reg  r_2725; // @[Reg.scala 16:16]
  reg  r_2726; // @[Reg.scala 16:16]
  reg  r_2727; // @[Reg.scala 16:16]
  reg  r_2728; // @[Reg.scala 16:16]
  reg  r_2729; // @[Reg.scala 16:16]
  reg  r_2730; // @[Reg.scala 16:16]
  reg  r_2731; // @[Reg.scala 16:16]
  reg  r_2732; // @[Reg.scala 16:16]
  reg  r_2733; // @[Reg.scala 16:16]
  reg  r_2734; // @[Reg.scala 16:16]
  reg  r_2735; // @[Reg.scala 16:16]
  reg  r_2736; // @[Reg.scala 16:16]
  reg  r_2737; // @[Reg.scala 16:16]
  reg  r_2738; // @[Reg.scala 16:16]
  reg  r_2739; // @[Reg.scala 16:16]
  reg  r_2740; // @[Reg.scala 16:16]
  reg  r_2741; // @[Reg.scala 16:16]
  reg  r_2742; // @[Reg.scala 16:16]
  reg  r_2743; // @[Reg.scala 16:16]
  reg  r_2744; // @[Reg.scala 16:16]
  reg  r_2745; // @[Reg.scala 16:16]
  reg  r_2746; // @[Reg.scala 16:16]
  reg  r_2747; // @[Reg.scala 16:16]
  reg  r_2748; // @[Reg.scala 16:16]
  reg  r_2749; // @[Reg.scala 16:16]
  reg  r_2750; // @[Reg.scala 16:16]
  reg  r_2751; // @[Reg.scala 16:16]
  reg  r_2752; // @[Reg.scala 16:16]
  reg  r_2753; // @[Reg.scala 16:16]
  reg  r_2754; // @[Reg.scala 16:16]
  reg  r_2755; // @[Reg.scala 16:16]
  reg  r_2756; // @[Reg.scala 16:16]
  reg  r_2757; // @[Reg.scala 16:16]
  reg  r_2758; // @[Reg.scala 16:16]
  reg  r_2759; // @[Reg.scala 16:16]
  reg  r_2760; // @[Reg.scala 16:16]
  reg  r_2761; // @[Reg.scala 16:16]
  reg  r_2762; // @[Reg.scala 16:16]
  reg  r_2763; // @[Reg.scala 16:16]
  reg  r_2764; // @[Reg.scala 16:16]
  reg  r_2765; // @[Reg.scala 16:16]
  reg  r_2766; // @[Reg.scala 16:16]
  reg  r_2767; // @[Reg.scala 16:16]
  reg  r_2768; // @[Reg.scala 16:16]
  reg  r_2769; // @[Reg.scala 16:16]
  reg  r_2770; // @[Reg.scala 16:16]
  reg  r_2771; // @[Reg.scala 16:16]
  reg  r_2772; // @[Reg.scala 16:16]
  reg  r_2773; // @[Reg.scala 16:16]
  reg  r_2774; // @[Reg.scala 16:16]
  reg  r_2775; // @[Reg.scala 16:16]
  reg  r_2776; // @[Reg.scala 16:16]
  reg  r_2777; // @[Reg.scala 16:16]
  reg  r_2778; // @[Reg.scala 16:16]
  reg  r_2779; // @[Reg.scala 16:16]
  reg  r_2780; // @[Reg.scala 16:16]
  reg  r_2781; // @[Reg.scala 16:16]
  reg  r_2782; // @[Reg.scala 16:16]
  reg  r_2783; // @[Reg.scala 16:16]
  reg  r_2784; // @[Reg.scala 16:16]
  reg  r_2785; // @[Reg.scala 16:16]
  reg  r_2786; // @[Reg.scala 16:16]
  reg  r_2787; // @[Reg.scala 16:16]
  reg  r_2788; // @[Reg.scala 16:16]
  reg  r_2789; // @[Reg.scala 16:16]
  reg  r_2790; // @[Reg.scala 16:16]
  reg  r_2791; // @[Reg.scala 16:16]
  reg  r_2792; // @[Reg.scala 16:16]
  reg  r_2793; // @[Reg.scala 16:16]
  reg  r_2794; // @[Reg.scala 16:16]
  reg  r_2795; // @[Reg.scala 16:16]
  reg  r_2796; // @[Reg.scala 16:16]
  reg  r_2797; // @[Reg.scala 16:16]
  reg  r_2798; // @[Reg.scala 16:16]
  reg  r_2799; // @[Reg.scala 16:16]
  reg  r_2800; // @[Reg.scala 16:16]
  reg  r_2801; // @[Reg.scala 16:16]
  reg  r_2802; // @[Reg.scala 16:16]
  reg  r_2803; // @[Reg.scala 16:16]
  reg  r_2804; // @[Reg.scala 16:16]
  reg  r_2805; // @[Reg.scala 16:16]
  reg  r_2806; // @[Reg.scala 16:16]
  reg  r_2807; // @[Reg.scala 16:16]
  reg  r_2808; // @[Reg.scala 16:16]
  reg  r_2809; // @[Reg.scala 16:16]
  reg  r_2810; // @[Reg.scala 16:16]
  reg  r_2811; // @[Reg.scala 16:16]
  reg  r_2812; // @[Reg.scala 16:16]
  reg  r_2813; // @[Reg.scala 16:16]
  reg  r_2814; // @[Reg.scala 16:16]
  reg  r_2815; // @[Reg.scala 16:16]
  reg  r_2816; // @[Reg.scala 16:16]
  reg  r_2817; // @[Reg.scala 16:16]
  reg  r_2818; // @[Reg.scala 16:16]
  reg  r_2819; // @[Reg.scala 16:16]
  reg  r_2820; // @[Reg.scala 16:16]
  reg  r_2821; // @[Reg.scala 16:16]
  reg  r_2822; // @[Reg.scala 16:16]
  reg  r_2823; // @[Reg.scala 16:16]
  reg  r_2824; // @[Reg.scala 16:16]
  reg  r_2825; // @[Reg.scala 16:16]
  reg  r_2826; // @[Reg.scala 16:16]
  reg  r_2827; // @[Reg.scala 16:16]
  reg  r_2828; // @[Reg.scala 16:16]
  reg  r_2829; // @[Reg.scala 16:16]
  reg  r_2830; // @[Reg.scala 16:16]
  reg  r_2831; // @[Reg.scala 16:16]
  reg  r_2832; // @[Reg.scala 16:16]
  reg  r_2833; // @[Reg.scala 16:16]
  reg  r_2834; // @[Reg.scala 16:16]
  reg  r_2835; // @[Reg.scala 16:16]
  reg  r_2836; // @[Reg.scala 16:16]
  reg  r_2837; // @[Reg.scala 16:16]
  reg  r_2838; // @[Reg.scala 16:16]
  reg  r_2839; // @[Reg.scala 16:16]
  reg  r_2840; // @[Reg.scala 16:16]
  reg  r_2841; // @[Reg.scala 16:16]
  reg  r_2842; // @[Reg.scala 16:16]
  reg  r_2843; // @[Reg.scala 16:16]
  reg  r_2844; // @[Reg.scala 16:16]
  reg  r_2845; // @[Reg.scala 16:16]
  reg  r_2846; // @[Reg.scala 16:16]
  reg  r_2847; // @[Reg.scala 16:16]
  reg  r_2848; // @[Reg.scala 16:16]
  reg  r_2849; // @[Reg.scala 16:16]
  reg  r_2850; // @[Reg.scala 16:16]
  reg  r_2851; // @[Reg.scala 16:16]
  reg  r_2852; // @[Reg.scala 16:16]
  reg  r_2853; // @[Reg.scala 16:16]
  reg  r_2854; // @[Reg.scala 16:16]
  reg  r_2855; // @[Reg.scala 16:16]
  reg  r_2856; // @[Reg.scala 16:16]
  reg  r_2857; // @[Reg.scala 16:16]
  reg  r_2858; // @[Reg.scala 16:16]
  reg  r_2859; // @[Reg.scala 16:16]
  reg  r_2860; // @[Reg.scala 16:16]
  reg  r_2861; // @[Reg.scala 16:16]
  reg  r_2862; // @[Reg.scala 16:16]
  reg  r_2863; // @[Reg.scala 16:16]
  reg  r_2864; // @[Reg.scala 16:16]
  reg  r_2865; // @[Reg.scala 16:16]
  reg  r_2866; // @[Reg.scala 16:16]
  reg  r_2867; // @[Reg.scala 16:16]
  reg  r_2868; // @[Reg.scala 16:16]
  reg  r_2869; // @[Reg.scala 16:16]
  reg  r_2870; // @[Reg.scala 16:16]
  wire  s_0_714 = m_2462_io_s; // @[MUL.scala 252:21]
  wire  c_0_714 = m_2462_io_cout; // @[MUL.scala 253:22]
  wire  s_0_715 = m_2463_io_s; // @[MUL.scala 252:21]
  wire  c_0_715 = m_2463_io_cout; // @[MUL.scala 253:22]
  wire  s_0_716 = m_2464_io_s; // @[MUL.scala 252:21]
  wire  c_0_716 = m_2464_io_cout; // @[MUL.scala 253:22]
  wire  s_0_717 = m_2465_io_s; // @[MUL.scala 252:21]
  wire  c_0_717 = m_2465_io_cout; // @[MUL.scala 253:22]
  wire  s_0_718 = m_2466_io_s; // @[MUL.scala 252:21]
  wire  c_0_718 = m_2466_io_cout; // @[MUL.scala 253:22]
  wire  s_0_719 = m_2467_io_s; // @[MUL.scala 252:21]
  wire  c_0_719 = m_2467_io_cout; // @[MUL.scala 253:22]
  wire  s_0_720 = m_2468_io_s; // @[MUL.scala 252:21]
  wire  c_0_720 = m_2468_io_cout; // @[MUL.scala 253:22]
  wire  s_0_721 = m_2469_io_s; // @[MUL.scala 252:21]
  wire  c_0_721 = m_2469_io_cout; // @[MUL.scala 253:22]
  wire  s_0_722 = m_2470_io_s; // @[MUL.scala 252:21]
  wire  c_0_722 = m_2470_io_cout; // @[MUL.scala 253:22]
  wire  s_0_723 = m_2471_io_s; // @[MUL.scala 252:21]
  wire  c_0_723 = m_2471_io_cout; // @[MUL.scala 253:22]
  wire  s_0_724 = m_2472_io_s; // @[MUL.scala 252:21]
  wire  c_0_724 = m_2472_io_cout; // @[MUL.scala 253:22]
  wire  s_0_725 = m_2473_io_s; // @[MUL.scala 252:21]
  wire  c_0_725 = m_2473_io_cout; // @[MUL.scala 253:22]
  wire  s_0_726 = m_2474_io_s; // @[MUL.scala 252:21]
  wire  c_0_726 = m_2474_io_cout; // @[MUL.scala 253:22]
  wire  s_0_727 = m_2475_io_s; // @[MUL.scala 252:21]
  wire  c_0_727 = m_2475_io_cout; // @[MUL.scala 253:22]
  wire  s_0_728 = m_2476_io_s; // @[MUL.scala 252:21]
  wire  c_0_728 = m_2476_io_cout; // @[MUL.scala 253:22]
  wire  s_0_729 = m_2477_io_s; // @[MUL.scala 252:21]
  wire  c_0_729 = m_2477_io_cout; // @[MUL.scala 253:22]
  wire  s_0_730 = m_2478_io_s; // @[MUL.scala 252:21]
  wire  c_0_730 = m_2478_io_cout; // @[MUL.scala 253:22]
  wire  s_0_731 = m_2479_io_s; // @[MUL.scala 252:21]
  wire  c_0_731 = m_2479_io_cout; // @[MUL.scala 253:22]
  wire  s_0_732 = m_2480_io_s; // @[MUL.scala 252:21]
  wire  c_0_732 = m_2480_io_cout; // @[MUL.scala 253:22]
  wire  s_0_733 = m_2481_io_s; // @[MUL.scala 252:21]
  wire  c_0_733 = m_2481_io_cout; // @[MUL.scala 253:22]
  wire  s_0_734 = m_2482_io_s; // @[MUL.scala 252:21]
  wire  c_0_734 = m_2482_io_cout; // @[MUL.scala 253:22]
  wire [7:0] sum_lo_lo_lo_lo = {m_2411_io_out_0,m_2286_io_out_0,m_2139_io_out_0,m_1954_io_out_0,r_2311,r_2310,r_2309,
    r_2308}; // @[Cat.scala 31:58]
  wire [15:0] sum_lo_lo_lo = {m_2419_io_out_0,m_2418_io_out_0,m_2417_io_out_0,m_2416_io_out_0,m_2415_io_out_0,
    m_2414_io_out_0,m_2413_io_out_0,m_2412_io_out_0,sum_lo_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] sum_lo_lo_hi_lo = {m_2427_io_out_0,m_2426_io_out_0,m_2425_io_out_0,m_2424_io_out_0,m_2423_io_out_0,
    m_2422_io_out_0,m_2421_io_out_0,m_2420_io_out_0}; // @[Cat.scala 31:58]
  wire [31:0] sum_lo_lo = {m_2435_io_out_0,m_2434_io_out_0,m_2433_io_out_0,m_2432_io_out_0,m_2431_io_out_0,
    m_2430_io_out_0,m_2429_io_out_0,m_2428_io_out_0,sum_lo_lo_hi_lo,sum_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] sum_lo_hi_lo_lo = {m_2443_io_out_0,m_2442_io_out_0,m_2441_io_out_0,m_2440_io_out_0,m_2439_io_out_0,
    m_2438_io_out_0,m_2437_io_out_0,m_2436_io_out_0}; // @[Cat.scala 31:58]
  wire [7:0] sum_lo_hi_hi_lo = {m_2459_io_out_0,m_2458_io_out_0,m_2457_io_out_0,m_2456_io_out_0,m_2455_io_out_0,
    m_2454_io_out_0,m_2453_io_out_0,m_2452_io_out_0}; // @[Cat.scala 31:58]
  wire [16:0] sum_lo_hi_hi = {s_0_720,s_0_719,s_0_718,s_0_717,s_0_716,s_0_715,s_0_714,m_2461_io_out_0,m_2460_io_out_0,
    sum_lo_hi_hi_lo}; // @[Cat.scala 31:58]
  wire [32:0] sum_lo_hi = {sum_lo_hi_hi,m_2451_io_out_0,m_2450_io_out_0,m_2449_io_out_0,m_2448_io_out_0,m_2447_io_out_0,
    m_2446_io_out_0,m_2445_io_out_0,m_2444_io_out_0,sum_lo_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] sum_hi_lo_lo_lo = {s_0_728,s_0_727,s_0_726,s_0_725,s_0_724,s_0_723,s_0_722,s_0_721}; // @[Cat.scala 31:58]
  wire [7:0] sum_hi_lo_hi_lo = {m_2492_io_out_0,m_2491_io_out_0,m_2490_io_out_0,m_2489_io_out_0,m_2488_io_out_0,
    m_2487_io_out_0,m_2486_io_out_0,m_2485_io_out_0}; // @[Cat.scala 31:58]
  wire [16:0] sum_hi_lo_hi = {m_2501_io_out_0,m_2500_io_out_0,m_2499_io_out_0,m_2498_io_out_0,m_2497_io_out_0,
    m_2496_io_out_0,m_2495_io_out_0,m_2494_io_out_0,m_2493_io_out_0,sum_hi_lo_hi_lo}; // @[Cat.scala 31:58]
  wire [32:0] sum_hi_lo = {sum_hi_lo_hi,m_2484_io_out_0,m_2483_io_out_0,s_0_734,s_0_733,s_0_732,s_0_731,s_0_730,s_0_729,
    sum_hi_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] sum_hi_hi_lo_lo = {m_2509_io_out_0,m_2508_io_out_0,m_2507_io_out_0,m_2506_io_out_0,m_2505_io_out_0,
    m_2504_io_out_0,m_2503_io_out_0,m_2502_io_out_0}; // @[Cat.scala 31:58]
  wire [7:0] sum_hi_hi_hi_lo = {m_2525_io_out_0,m_2524_io_out_0,m_2523_io_out_0,m_2522_io_out_0,m_2521_io_out_0,
    m_2520_io_out_0,m_2519_io_out_0,m_2518_io_out_0}; // @[Cat.scala 31:58]
  wire [16:0] sum_hi_hi_hi = {m_2534_io_out_0,m_2533_io_out_0,m_2532_io_out_0,m_2531_io_out_0,m_2530_io_out_0,
    m_2529_io_out_0,m_2528_io_out_0,m_2527_io_out_0,m_2526_io_out_0,sum_hi_hi_hi_lo}; // @[Cat.scala 31:58]
  wire [32:0] sum_hi_hi = {sum_hi_hi_hi,m_2517_io_out_0,m_2516_io_out_0,m_2515_io_out_0,m_2514_io_out_0,m_2513_io_out_0,
    m_2512_io_out_0,m_2511_io_out_0,m_2510_io_out_0,sum_hi_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [130:0] sum = {sum_hi_hi,sum_hi_lo,sum_lo_hi,sum_lo_lo}; // @[Cat.scala 31:58]
  wire [6:0] carry_lo_lo_lo_lo = {m_2417_io_out_1,m_2416_io_out_1,m_2415_io_out_1,m_2414_io_out_1,m_2413_io_out_1,
    m_2412_io_out_1,m_2411_io_out_1}; // @[Cat.scala 31:58]
  wire [14:0] carry_lo_lo_lo = {m_2425_io_out_1,m_2424_io_out_1,m_2423_io_out_1,m_2422_io_out_1,m_2421_io_out_1,
    m_2420_io_out_1,m_2419_io_out_1,m_2418_io_out_1,carry_lo_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [6:0] carry_lo_lo_hi_lo = {m_2432_io_out_1,m_2431_io_out_1,m_2430_io_out_1,m_2429_io_out_1,m_2428_io_out_1,
    m_2427_io_out_1,m_2426_io_out_1}; // @[Cat.scala 31:58]
  wire [29:0] carry_lo_lo = {m_2440_io_out_1,m_2439_io_out_1,m_2438_io_out_1,m_2437_io_out_1,m_2436_io_out_1,
    m_2435_io_out_1,m_2434_io_out_1,m_2433_io_out_1,carry_lo_lo_hi_lo,carry_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [6:0] carry_lo_hi_lo_lo = {m_2447_io_out_1,m_2446_io_out_1,m_2445_io_out_1,m_2444_io_out_1,m_2443_io_out_1,
    m_2442_io_out_1,m_2441_io_out_1}; // @[Cat.scala 31:58]
  wire [14:0] carry_lo_hi_lo = {m_2455_io_out_1,m_2454_io_out_1,m_2453_io_out_1,m_2452_io_out_1,m_2451_io_out_1,
    m_2450_io_out_1,m_2449_io_out_1,m_2448_io_out_1,carry_lo_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] carry_lo_hi_hi_lo = {c_0_715,c_0_714,m_2461_io_out_1,m_2460_io_out_1,m_2459_io_out_1,m_2458_io_out_1,
    m_2457_io_out_1,m_2456_io_out_1}; // @[Cat.scala 31:58]
  wire [30:0] carry_lo_hi = {c_0_723,c_0_722,c_0_721,c_0_720,c_0_719,c_0_718,c_0_717,c_0_716,carry_lo_hi_hi_lo,
    carry_lo_hi_lo}; // @[Cat.scala 31:58]
  wire [6:0] carry_hi_lo_lo_lo = {c_0_730,c_0_729,c_0_728,c_0_727,c_0_726,c_0_725,c_0_724}; // @[Cat.scala 31:58]
  wire [14:0] carry_hi_lo_lo = {m_2486_io_out_1,m_2485_io_out_1,m_2484_io_out_1,m_2483_io_out_1,c_0_734,c_0_733,c_0_732,
    c_0_731,carry_hi_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] carry_hi_lo_hi_lo = {m_2494_io_out_1,m_2493_io_out_1,m_2492_io_out_1,m_2491_io_out_1,m_2490_io_out_1,
    m_2489_io_out_1,m_2488_io_out_1,m_2487_io_out_1}; // @[Cat.scala 31:58]
  wire [30:0] carry_hi_lo = {m_2502_io_out_1,m_2501_io_out_1,m_2500_io_out_1,m_2499_io_out_1,m_2498_io_out_1,
    m_2497_io_out_1,m_2496_io_out_1,m_2495_io_out_1,carry_hi_lo_hi_lo,carry_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [6:0] carry_hi_hi_lo_lo = {m_2509_io_out_1,m_2508_io_out_1,m_2507_io_out_1,m_2506_io_out_1,m_2505_io_out_1,
    m_2504_io_out_1,m_2503_io_out_1}; // @[Cat.scala 31:58]
  wire [14:0] carry_hi_hi_lo = {m_2517_io_out_1,m_2516_io_out_1,m_2515_io_out_1,m_2514_io_out_1,m_2513_io_out_1,
    m_2512_io_out_1,m_2511_io_out_1,m_2510_io_out_1,carry_hi_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] carry_hi_hi_hi_lo = {m_2525_io_out_1,m_2524_io_out_1,m_2523_io_out_1,m_2522_io_out_1,m_2521_io_out_1,
    m_2520_io_out_1,m_2519_io_out_1,m_2518_io_out_1}; // @[Cat.scala 31:58]
  wire [30:0] carry_hi_hi = {m_2533_io_out_1,m_2532_io_out_1,m_2531_io_out_1,m_2530_io_out_1,m_2529_io_out_1,
    m_2528_io_out_1,m_2527_io_out_1,m_2526_io_out_1,carry_hi_hi_hi_lo,carry_hi_hi_lo}; // @[Cat.scala 31:58]
  wire [130:0] cout = {carry_hi_hi,carry_hi_lo,carry_lo_hi,carry_lo_lo,8'h0}; // @[Cat.scala 31:58]
  wire [130:0] result = sum + cout; // @[MUL.scala 332:20]
  reg [7:0] count; // @[MUL.scala 334:22]
  wire [7:0] _count_T_5 = count + 8'h1; // @[MUL.scala 336:81]
  Improved_Partial_product m ( // @[MUL.scala 81:21]
    .io_y_3(m_io_y_3),
    .io_x(m_io_x),
    .io_p(m_io_p),
    .io_carry(m_io_carry)
  );
  Improved_Partial_product m_1 ( // @[MUL.scala 81:21]
    .io_y_3(m_1_io_y_3),
    .io_x(m_1_io_x),
    .io_p(m_1_io_p),
    .io_carry(m_1_io_carry)
  );
  Improved_Partial_product m_2 ( // @[MUL.scala 81:21]
    .io_y_3(m_2_io_y_3),
    .io_x(m_2_io_x),
    .io_p(m_2_io_p),
    .io_carry(m_2_io_carry)
  );
  Improved_Partial_product m_3 ( // @[MUL.scala 81:21]
    .io_y_3(m_3_io_y_3),
    .io_x(m_3_io_x),
    .io_p(m_3_io_p),
    .io_carry(m_3_io_carry)
  );
  Improved_Partial_product m_4 ( // @[MUL.scala 81:21]
    .io_y_3(m_4_io_y_3),
    .io_x(m_4_io_x),
    .io_p(m_4_io_p),
    .io_carry(m_4_io_carry)
  );
  Improved_Partial_product m_5 ( // @[MUL.scala 81:21]
    .io_y_3(m_5_io_y_3),
    .io_x(m_5_io_x),
    .io_p(m_5_io_p),
    .io_carry(m_5_io_carry)
  );
  Improved_Partial_product m_6 ( // @[MUL.scala 81:21]
    .io_y_3(m_6_io_y_3),
    .io_x(m_6_io_x),
    .io_p(m_6_io_p),
    .io_carry(m_6_io_carry)
  );
  Improved_Partial_product m_7 ( // @[MUL.scala 81:21]
    .io_y_3(m_7_io_y_3),
    .io_x(m_7_io_x),
    .io_p(m_7_io_p),
    .io_carry(m_7_io_carry)
  );
  Improved_Partial_product m_8 ( // @[MUL.scala 81:21]
    .io_y_3(m_8_io_y_3),
    .io_x(m_8_io_x),
    .io_p(m_8_io_p),
    .io_carry(m_8_io_carry)
  );
  Improved_Partial_product m_9 ( // @[MUL.scala 81:21]
    .io_y_3(m_9_io_y_3),
    .io_x(m_9_io_x),
    .io_p(m_9_io_p),
    .io_carry(m_9_io_carry)
  );
  Improved_Partial_product m_10 ( // @[MUL.scala 81:21]
    .io_y_3(m_10_io_y_3),
    .io_x(m_10_io_x),
    .io_p(m_10_io_p),
    .io_carry(m_10_io_carry)
  );
  Improved_Partial_product m_11 ( // @[MUL.scala 81:21]
    .io_y_3(m_11_io_y_3),
    .io_x(m_11_io_x),
    .io_p(m_11_io_p),
    .io_carry(m_11_io_carry)
  );
  Improved_Partial_product m_12 ( // @[MUL.scala 81:21]
    .io_y_3(m_12_io_y_3),
    .io_x(m_12_io_x),
    .io_p(m_12_io_p),
    .io_carry(m_12_io_carry)
  );
  Improved_Partial_product m_13 ( // @[MUL.scala 81:21]
    .io_y_3(m_13_io_y_3),
    .io_x(m_13_io_x),
    .io_p(m_13_io_p),
    .io_carry(m_13_io_carry)
  );
  Improved_Partial_product m_14 ( // @[MUL.scala 81:21]
    .io_y_3(m_14_io_y_3),
    .io_x(m_14_io_x),
    .io_p(m_14_io_p),
    .io_carry(m_14_io_carry)
  );
  Improved_Partial_product m_15 ( // @[MUL.scala 81:21]
    .io_y_3(m_15_io_y_3),
    .io_x(m_15_io_x),
    .io_p(m_15_io_p),
    .io_carry(m_15_io_carry)
  );
  Improved_Partial_product m_16 ( // @[MUL.scala 81:21]
    .io_y_3(m_16_io_y_3),
    .io_x(m_16_io_x),
    .io_p(m_16_io_p),
    .io_carry(m_16_io_carry)
  );
  Improved_Partial_product m_17 ( // @[MUL.scala 81:21]
    .io_y_3(m_17_io_y_3),
    .io_x(m_17_io_x),
    .io_p(m_17_io_p),
    .io_carry(m_17_io_carry)
  );
  Improved_Partial_product m_18 ( // @[MUL.scala 81:21]
    .io_y_3(m_18_io_y_3),
    .io_x(m_18_io_x),
    .io_p(m_18_io_p),
    .io_carry(m_18_io_carry)
  );
  Improved_Partial_product m_19 ( // @[MUL.scala 81:21]
    .io_y_3(m_19_io_y_3),
    .io_x(m_19_io_x),
    .io_p(m_19_io_p),
    .io_carry(m_19_io_carry)
  );
  Improved_Partial_product m_20 ( // @[MUL.scala 81:21]
    .io_y_3(m_20_io_y_3),
    .io_x(m_20_io_x),
    .io_p(m_20_io_p),
    .io_carry(m_20_io_carry)
  );
  Improved_Partial_product m_21 ( // @[MUL.scala 81:21]
    .io_y_3(m_21_io_y_3),
    .io_x(m_21_io_x),
    .io_p(m_21_io_p),
    .io_carry(m_21_io_carry)
  );
  Improved_Partial_product m_22 ( // @[MUL.scala 81:21]
    .io_y_3(m_22_io_y_3),
    .io_x(m_22_io_x),
    .io_p(m_22_io_p),
    .io_carry(m_22_io_carry)
  );
  Improved_Partial_product m_23 ( // @[MUL.scala 81:21]
    .io_y_3(m_23_io_y_3),
    .io_x(m_23_io_x),
    .io_p(m_23_io_p),
    .io_carry(m_23_io_carry)
  );
  Improved_Partial_product m_24 ( // @[MUL.scala 81:21]
    .io_y_3(m_24_io_y_3),
    .io_x(m_24_io_x),
    .io_p(m_24_io_p),
    .io_carry(m_24_io_carry)
  );
  Improved_Partial_product m_25 ( // @[MUL.scala 81:21]
    .io_y_3(m_25_io_y_3),
    .io_x(m_25_io_x),
    .io_p(m_25_io_p),
    .io_carry(m_25_io_carry)
  );
  Improved_Partial_product m_26 ( // @[MUL.scala 81:21]
    .io_y_3(m_26_io_y_3),
    .io_x(m_26_io_x),
    .io_p(m_26_io_p),
    .io_carry(m_26_io_carry)
  );
  Improved_Partial_product m_27 ( // @[MUL.scala 81:21]
    .io_y_3(m_27_io_y_3),
    .io_x(m_27_io_x),
    .io_p(m_27_io_p),
    .io_carry(m_27_io_carry)
  );
  Improved_Partial_product m_28 ( // @[MUL.scala 81:21]
    .io_y_3(m_28_io_y_3),
    .io_x(m_28_io_x),
    .io_p(m_28_io_p),
    .io_carry(m_28_io_carry)
  );
  Improved_Partial_product m_29 ( // @[MUL.scala 81:21]
    .io_y_3(m_29_io_y_3),
    .io_x(m_29_io_x),
    .io_p(m_29_io_p),
    .io_carry(m_29_io_carry)
  );
  Improved_Partial_product m_30 ( // @[MUL.scala 81:21]
    .io_y_3(m_30_io_y_3),
    .io_x(m_30_io_x),
    .io_p(m_30_io_p),
    .io_carry(m_30_io_carry)
  );
  Improved_Partial_product m_31 ( // @[MUL.scala 81:21]
    .io_y_3(m_31_io_y_3),
    .io_x(m_31_io_x),
    .io_p(m_31_io_p),
    .io_carry(m_31_io_carry)
  );
  Improved_Partial_product m_32 ( // @[MUL.scala 81:21]
    .io_y_3(m_32_io_y_3),
    .io_x(m_32_io_x),
    .io_p(m_32_io_p),
    .io_carry(m_32_io_carry)
  );
  Half_Adder m_33 ( // @[MUL.scala 124:19]
    .io_in_0(m_33_io_in_0),
    .io_in_1(m_33_io_in_1),
    .io_out_0(m_33_io_out_0),
    .io_out_1(m_33_io_out_1)
  );
  Half_Adder m_34 ( // @[MUL.scala 124:19]
    .io_in_0(m_34_io_in_0),
    .io_in_1(m_34_io_in_1),
    .io_out_0(m_34_io_out_0),
    .io_out_1(m_34_io_out_1)
  );
  Adder m_35 ( // @[MUL.scala 102:19]
    .io_x1(m_35_io_x1),
    .io_x2(m_35_io_x2),
    .io_x3(m_35_io_x3),
    .io_s(m_35_io_s),
    .io_cout(m_35_io_cout)
  );
  Adder m_36 ( // @[MUL.scala 102:19]
    .io_x1(m_36_io_x1),
    .io_x2(m_36_io_x2),
    .io_x3(m_36_io_x3),
    .io_s(m_36_io_s),
    .io_cout(m_36_io_cout)
  );
  Adder m_37 ( // @[MUL.scala 102:19]
    .io_x1(m_37_io_x1),
    .io_x2(m_37_io_x2),
    .io_x3(m_37_io_x3),
    .io_s(m_37_io_s),
    .io_cout(m_37_io_cout)
  );
  Adder m_38 ( // @[MUL.scala 102:19]
    .io_x1(m_38_io_x1),
    .io_x2(m_38_io_x2),
    .io_x3(m_38_io_x3),
    .io_s(m_38_io_s),
    .io_cout(m_38_io_cout)
  );
  Adder m_39 ( // @[MUL.scala 102:19]
    .io_x1(m_39_io_x1),
    .io_x2(m_39_io_x2),
    .io_x3(m_39_io_x3),
    .io_s(m_39_io_s),
    .io_cout(m_39_io_cout)
  );
  Half_Adder m_40 ( // @[MUL.scala 124:19]
    .io_in_0(m_40_io_in_0),
    .io_in_1(m_40_io_in_1),
    .io_out_0(m_40_io_out_0),
    .io_out_1(m_40_io_out_1)
  );
  Adder m_41 ( // @[MUL.scala 102:19]
    .io_x1(m_41_io_x1),
    .io_x2(m_41_io_x2),
    .io_x3(m_41_io_x3),
    .io_s(m_41_io_s),
    .io_cout(m_41_io_cout)
  );
  Half_Adder m_42 ( // @[MUL.scala 124:19]
    .io_in_0(m_42_io_in_0),
    .io_in_1(m_42_io_in_1),
    .io_out_0(m_42_io_out_0),
    .io_out_1(m_42_io_out_1)
  );
  Adder m_43 ( // @[MUL.scala 102:19]
    .io_x1(m_43_io_x1),
    .io_x2(m_43_io_x2),
    .io_x3(m_43_io_x3),
    .io_s(m_43_io_s),
    .io_cout(m_43_io_cout)
  );
  Adder m_44 ( // @[MUL.scala 102:19]
    .io_x1(m_44_io_x1),
    .io_x2(m_44_io_x2),
    .io_x3(m_44_io_x3),
    .io_s(m_44_io_s),
    .io_cout(m_44_io_cout)
  );
  Adder m_45 ( // @[MUL.scala 102:19]
    .io_x1(m_45_io_x1),
    .io_x2(m_45_io_x2),
    .io_x3(m_45_io_x3),
    .io_s(m_45_io_s),
    .io_cout(m_45_io_cout)
  );
  Adder m_46 ( // @[MUL.scala 102:19]
    .io_x1(m_46_io_x1),
    .io_x2(m_46_io_x2),
    .io_x3(m_46_io_x3),
    .io_s(m_46_io_s),
    .io_cout(m_46_io_cout)
  );
  Adder m_47 ( // @[MUL.scala 102:19]
    .io_x1(m_47_io_x1),
    .io_x2(m_47_io_x2),
    .io_x3(m_47_io_x3),
    .io_s(m_47_io_s),
    .io_cout(m_47_io_cout)
  );
  Adder m_48 ( // @[MUL.scala 102:19]
    .io_x1(m_48_io_x1),
    .io_x2(m_48_io_x2),
    .io_x3(m_48_io_x3),
    .io_s(m_48_io_s),
    .io_cout(m_48_io_cout)
  );
  Adder m_49 ( // @[MUL.scala 102:19]
    .io_x1(m_49_io_x1),
    .io_x2(m_49_io_x2),
    .io_x3(m_49_io_x3),
    .io_s(m_49_io_s),
    .io_cout(m_49_io_cout)
  );
  Adder m_50 ( // @[MUL.scala 102:19]
    .io_x1(m_50_io_x1),
    .io_x2(m_50_io_x2),
    .io_x3(m_50_io_x3),
    .io_s(m_50_io_s),
    .io_cout(m_50_io_cout)
  );
  Adder m_51 ( // @[MUL.scala 102:19]
    .io_x1(m_51_io_x1),
    .io_x2(m_51_io_x2),
    .io_x3(m_51_io_x3),
    .io_s(m_51_io_s),
    .io_cout(m_51_io_cout)
  );
  Adder m_52 ( // @[MUL.scala 102:19]
    .io_x1(m_52_io_x1),
    .io_x2(m_52_io_x2),
    .io_x3(m_52_io_x3),
    .io_s(m_52_io_s),
    .io_cout(m_52_io_cout)
  );
  Half_Adder m_53 ( // @[MUL.scala 124:19]
    .io_in_0(m_53_io_in_0),
    .io_in_1(m_53_io_in_1),
    .io_out_0(m_53_io_out_0),
    .io_out_1(m_53_io_out_1)
  );
  Adder m_54 ( // @[MUL.scala 102:19]
    .io_x1(m_54_io_x1),
    .io_x2(m_54_io_x2),
    .io_x3(m_54_io_x3),
    .io_s(m_54_io_s),
    .io_cout(m_54_io_cout)
  );
  Adder m_55 ( // @[MUL.scala 102:19]
    .io_x1(m_55_io_x1),
    .io_x2(m_55_io_x2),
    .io_x3(m_55_io_x3),
    .io_s(m_55_io_s),
    .io_cout(m_55_io_cout)
  );
  Half_Adder m_56 ( // @[MUL.scala 124:19]
    .io_in_0(m_56_io_in_0),
    .io_in_1(m_56_io_in_1),
    .io_out_0(m_56_io_out_0),
    .io_out_1(m_56_io_out_1)
  );
  Adder m_57 ( // @[MUL.scala 102:19]
    .io_x1(m_57_io_x1),
    .io_x2(m_57_io_x2),
    .io_x3(m_57_io_x3),
    .io_s(m_57_io_s),
    .io_cout(m_57_io_cout)
  );
  Adder m_58 ( // @[MUL.scala 102:19]
    .io_x1(m_58_io_x1),
    .io_x2(m_58_io_x2),
    .io_x3(m_58_io_x3),
    .io_s(m_58_io_s),
    .io_cout(m_58_io_cout)
  );
  Adder m_59 ( // @[MUL.scala 102:19]
    .io_x1(m_59_io_x1),
    .io_x2(m_59_io_x2),
    .io_x3(m_59_io_x3),
    .io_s(m_59_io_s),
    .io_cout(m_59_io_cout)
  );
  Adder m_60 ( // @[MUL.scala 102:19]
    .io_x1(m_60_io_x1),
    .io_x2(m_60_io_x2),
    .io_x3(m_60_io_x3),
    .io_s(m_60_io_s),
    .io_cout(m_60_io_cout)
  );
  Adder m_61 ( // @[MUL.scala 102:19]
    .io_x1(m_61_io_x1),
    .io_x2(m_61_io_x2),
    .io_x3(m_61_io_x3),
    .io_s(m_61_io_s),
    .io_cout(m_61_io_cout)
  );
  Adder m_62 ( // @[MUL.scala 102:19]
    .io_x1(m_62_io_x1),
    .io_x2(m_62_io_x2),
    .io_x3(m_62_io_x3),
    .io_s(m_62_io_s),
    .io_cout(m_62_io_cout)
  );
  Adder m_63 ( // @[MUL.scala 102:19]
    .io_x1(m_63_io_x1),
    .io_x2(m_63_io_x2),
    .io_x3(m_63_io_x3),
    .io_s(m_63_io_s),
    .io_cout(m_63_io_cout)
  );
  Adder m_64 ( // @[MUL.scala 102:19]
    .io_x1(m_64_io_x1),
    .io_x2(m_64_io_x2),
    .io_x3(m_64_io_x3),
    .io_s(m_64_io_s),
    .io_cout(m_64_io_cout)
  );
  Adder m_65 ( // @[MUL.scala 102:19]
    .io_x1(m_65_io_x1),
    .io_x2(m_65_io_x2),
    .io_x3(m_65_io_x3),
    .io_s(m_65_io_s),
    .io_cout(m_65_io_cout)
  );
  Adder m_66 ( // @[MUL.scala 102:19]
    .io_x1(m_66_io_x1),
    .io_x2(m_66_io_x2),
    .io_x3(m_66_io_x3),
    .io_s(m_66_io_s),
    .io_cout(m_66_io_cout)
  );
  Adder m_67 ( // @[MUL.scala 102:19]
    .io_x1(m_67_io_x1),
    .io_x2(m_67_io_x2),
    .io_x3(m_67_io_x3),
    .io_s(m_67_io_s),
    .io_cout(m_67_io_cout)
  );
  Adder m_68 ( // @[MUL.scala 102:19]
    .io_x1(m_68_io_x1),
    .io_x2(m_68_io_x2),
    .io_x3(m_68_io_x3),
    .io_s(m_68_io_s),
    .io_cout(m_68_io_cout)
  );
  Adder m_69 ( // @[MUL.scala 102:19]
    .io_x1(m_69_io_x1),
    .io_x2(m_69_io_x2),
    .io_x3(m_69_io_x3),
    .io_s(m_69_io_s),
    .io_cout(m_69_io_cout)
  );
  Adder m_70 ( // @[MUL.scala 102:19]
    .io_x1(m_70_io_x1),
    .io_x2(m_70_io_x2),
    .io_x3(m_70_io_x3),
    .io_s(m_70_io_s),
    .io_cout(m_70_io_cout)
  );
  Adder m_71 ( // @[MUL.scala 102:19]
    .io_x1(m_71_io_x1),
    .io_x2(m_71_io_x2),
    .io_x3(m_71_io_x3),
    .io_s(m_71_io_s),
    .io_cout(m_71_io_cout)
  );
  Half_Adder m_72 ( // @[MUL.scala 124:19]
    .io_in_0(m_72_io_in_0),
    .io_in_1(m_72_io_in_1),
    .io_out_0(m_72_io_out_0),
    .io_out_1(m_72_io_out_1)
  );
  Adder m_73 ( // @[MUL.scala 102:19]
    .io_x1(m_73_io_x1),
    .io_x2(m_73_io_x2),
    .io_x3(m_73_io_x3),
    .io_s(m_73_io_s),
    .io_cout(m_73_io_cout)
  );
  Adder m_74 ( // @[MUL.scala 102:19]
    .io_x1(m_74_io_x1),
    .io_x2(m_74_io_x2),
    .io_x3(m_74_io_x3),
    .io_s(m_74_io_s),
    .io_cout(m_74_io_cout)
  );
  Adder m_75 ( // @[MUL.scala 102:19]
    .io_x1(m_75_io_x1),
    .io_x2(m_75_io_x2),
    .io_x3(m_75_io_x3),
    .io_s(m_75_io_s),
    .io_cout(m_75_io_cout)
  );
  Half_Adder m_76 ( // @[MUL.scala 124:19]
    .io_in_0(m_76_io_in_0),
    .io_in_1(m_76_io_in_1),
    .io_out_0(m_76_io_out_0),
    .io_out_1(m_76_io_out_1)
  );
  Adder m_77 ( // @[MUL.scala 102:19]
    .io_x1(m_77_io_x1),
    .io_x2(m_77_io_x2),
    .io_x3(m_77_io_x3),
    .io_s(m_77_io_s),
    .io_cout(m_77_io_cout)
  );
  Adder m_78 ( // @[MUL.scala 102:19]
    .io_x1(m_78_io_x1),
    .io_x2(m_78_io_x2),
    .io_x3(m_78_io_x3),
    .io_s(m_78_io_s),
    .io_cout(m_78_io_cout)
  );
  Adder m_79 ( // @[MUL.scala 102:19]
    .io_x1(m_79_io_x1),
    .io_x2(m_79_io_x2),
    .io_x3(m_79_io_x3),
    .io_s(m_79_io_s),
    .io_cout(m_79_io_cout)
  );
  Adder m_80 ( // @[MUL.scala 102:19]
    .io_x1(m_80_io_x1),
    .io_x2(m_80_io_x2),
    .io_x3(m_80_io_x3),
    .io_s(m_80_io_s),
    .io_cout(m_80_io_cout)
  );
  Adder m_81 ( // @[MUL.scala 102:19]
    .io_x1(m_81_io_x1),
    .io_x2(m_81_io_x2),
    .io_x3(m_81_io_x3),
    .io_s(m_81_io_s),
    .io_cout(m_81_io_cout)
  );
  Adder m_82 ( // @[MUL.scala 102:19]
    .io_x1(m_82_io_x1),
    .io_x2(m_82_io_x2),
    .io_x3(m_82_io_x3),
    .io_s(m_82_io_s),
    .io_cout(m_82_io_cout)
  );
  Adder m_83 ( // @[MUL.scala 102:19]
    .io_x1(m_83_io_x1),
    .io_x2(m_83_io_x2),
    .io_x3(m_83_io_x3),
    .io_s(m_83_io_s),
    .io_cout(m_83_io_cout)
  );
  Adder m_84 ( // @[MUL.scala 102:19]
    .io_x1(m_84_io_x1),
    .io_x2(m_84_io_x2),
    .io_x3(m_84_io_x3),
    .io_s(m_84_io_s),
    .io_cout(m_84_io_cout)
  );
  Adder m_85 ( // @[MUL.scala 102:19]
    .io_x1(m_85_io_x1),
    .io_x2(m_85_io_x2),
    .io_x3(m_85_io_x3),
    .io_s(m_85_io_s),
    .io_cout(m_85_io_cout)
  );
  Adder m_86 ( // @[MUL.scala 102:19]
    .io_x1(m_86_io_x1),
    .io_x2(m_86_io_x2),
    .io_x3(m_86_io_x3),
    .io_s(m_86_io_s),
    .io_cout(m_86_io_cout)
  );
  Adder m_87 ( // @[MUL.scala 102:19]
    .io_x1(m_87_io_x1),
    .io_x2(m_87_io_x2),
    .io_x3(m_87_io_x3),
    .io_s(m_87_io_s),
    .io_cout(m_87_io_cout)
  );
  Adder m_88 ( // @[MUL.scala 102:19]
    .io_x1(m_88_io_x1),
    .io_x2(m_88_io_x2),
    .io_x3(m_88_io_x3),
    .io_s(m_88_io_s),
    .io_cout(m_88_io_cout)
  );
  Adder m_89 ( // @[MUL.scala 102:19]
    .io_x1(m_89_io_x1),
    .io_x2(m_89_io_x2),
    .io_x3(m_89_io_x3),
    .io_s(m_89_io_s),
    .io_cout(m_89_io_cout)
  );
  Adder m_90 ( // @[MUL.scala 102:19]
    .io_x1(m_90_io_x1),
    .io_x2(m_90_io_x2),
    .io_x3(m_90_io_x3),
    .io_s(m_90_io_s),
    .io_cout(m_90_io_cout)
  );
  Adder m_91 ( // @[MUL.scala 102:19]
    .io_x1(m_91_io_x1),
    .io_x2(m_91_io_x2),
    .io_x3(m_91_io_x3),
    .io_s(m_91_io_s),
    .io_cout(m_91_io_cout)
  );
  Adder m_92 ( // @[MUL.scala 102:19]
    .io_x1(m_92_io_x1),
    .io_x2(m_92_io_x2),
    .io_x3(m_92_io_x3),
    .io_s(m_92_io_s),
    .io_cout(m_92_io_cout)
  );
  Adder m_93 ( // @[MUL.scala 102:19]
    .io_x1(m_93_io_x1),
    .io_x2(m_93_io_x2),
    .io_x3(m_93_io_x3),
    .io_s(m_93_io_s),
    .io_cout(m_93_io_cout)
  );
  Adder m_94 ( // @[MUL.scala 102:19]
    .io_x1(m_94_io_x1),
    .io_x2(m_94_io_x2),
    .io_x3(m_94_io_x3),
    .io_s(m_94_io_s),
    .io_cout(m_94_io_cout)
  );
  Adder m_95 ( // @[MUL.scala 102:19]
    .io_x1(m_95_io_x1),
    .io_x2(m_95_io_x2),
    .io_x3(m_95_io_x3),
    .io_s(m_95_io_s),
    .io_cout(m_95_io_cout)
  );
  Adder m_96 ( // @[MUL.scala 102:19]
    .io_x1(m_96_io_x1),
    .io_x2(m_96_io_x2),
    .io_x3(m_96_io_x3),
    .io_s(m_96_io_s),
    .io_cout(m_96_io_cout)
  );
  Half_Adder m_97 ( // @[MUL.scala 124:19]
    .io_in_0(m_97_io_in_0),
    .io_in_1(m_97_io_in_1),
    .io_out_0(m_97_io_out_0),
    .io_out_1(m_97_io_out_1)
  );
  Adder m_98 ( // @[MUL.scala 102:19]
    .io_x1(m_98_io_x1),
    .io_x2(m_98_io_x2),
    .io_x3(m_98_io_x3),
    .io_s(m_98_io_s),
    .io_cout(m_98_io_cout)
  );
  Adder m_99 ( // @[MUL.scala 102:19]
    .io_x1(m_99_io_x1),
    .io_x2(m_99_io_x2),
    .io_x3(m_99_io_x3),
    .io_s(m_99_io_s),
    .io_cout(m_99_io_cout)
  );
  Adder m_100 ( // @[MUL.scala 102:19]
    .io_x1(m_100_io_x1),
    .io_x2(m_100_io_x2),
    .io_x3(m_100_io_x3),
    .io_s(m_100_io_s),
    .io_cout(m_100_io_cout)
  );
  Adder m_101 ( // @[MUL.scala 102:19]
    .io_x1(m_101_io_x1),
    .io_x2(m_101_io_x2),
    .io_x3(m_101_io_x3),
    .io_s(m_101_io_s),
    .io_cout(m_101_io_cout)
  );
  Half_Adder m_102 ( // @[MUL.scala 124:19]
    .io_in_0(m_102_io_in_0),
    .io_in_1(m_102_io_in_1),
    .io_out_0(m_102_io_out_0),
    .io_out_1(m_102_io_out_1)
  );
  Adder m_103 ( // @[MUL.scala 102:19]
    .io_x1(m_103_io_x1),
    .io_x2(m_103_io_x2),
    .io_x3(m_103_io_x3),
    .io_s(m_103_io_s),
    .io_cout(m_103_io_cout)
  );
  Adder m_104 ( // @[MUL.scala 102:19]
    .io_x1(m_104_io_x1),
    .io_x2(m_104_io_x2),
    .io_x3(m_104_io_x3),
    .io_s(m_104_io_s),
    .io_cout(m_104_io_cout)
  );
  Adder m_105 ( // @[MUL.scala 102:19]
    .io_x1(m_105_io_x1),
    .io_x2(m_105_io_x2),
    .io_x3(m_105_io_x3),
    .io_s(m_105_io_s),
    .io_cout(m_105_io_cout)
  );
  Adder m_106 ( // @[MUL.scala 102:19]
    .io_x1(m_106_io_x1),
    .io_x2(m_106_io_x2),
    .io_x3(m_106_io_x3),
    .io_s(m_106_io_s),
    .io_cout(m_106_io_cout)
  );
  Adder m_107 ( // @[MUL.scala 102:19]
    .io_x1(m_107_io_x1),
    .io_x2(m_107_io_x2),
    .io_x3(m_107_io_x3),
    .io_s(m_107_io_s),
    .io_cout(m_107_io_cout)
  );
  Adder m_108 ( // @[MUL.scala 102:19]
    .io_x1(m_108_io_x1),
    .io_x2(m_108_io_x2),
    .io_x3(m_108_io_x3),
    .io_s(m_108_io_s),
    .io_cout(m_108_io_cout)
  );
  Adder m_109 ( // @[MUL.scala 102:19]
    .io_x1(m_109_io_x1),
    .io_x2(m_109_io_x2),
    .io_x3(m_109_io_x3),
    .io_s(m_109_io_s),
    .io_cout(m_109_io_cout)
  );
  Adder m_110 ( // @[MUL.scala 102:19]
    .io_x1(m_110_io_x1),
    .io_x2(m_110_io_x2),
    .io_x3(m_110_io_x3),
    .io_s(m_110_io_s),
    .io_cout(m_110_io_cout)
  );
  Adder m_111 ( // @[MUL.scala 102:19]
    .io_x1(m_111_io_x1),
    .io_x2(m_111_io_x2),
    .io_x3(m_111_io_x3),
    .io_s(m_111_io_s),
    .io_cout(m_111_io_cout)
  );
  Adder m_112 ( // @[MUL.scala 102:19]
    .io_x1(m_112_io_x1),
    .io_x2(m_112_io_x2),
    .io_x3(m_112_io_x3),
    .io_s(m_112_io_s),
    .io_cout(m_112_io_cout)
  );
  Adder m_113 ( // @[MUL.scala 102:19]
    .io_x1(m_113_io_x1),
    .io_x2(m_113_io_x2),
    .io_x3(m_113_io_x3),
    .io_s(m_113_io_s),
    .io_cout(m_113_io_cout)
  );
  Adder m_114 ( // @[MUL.scala 102:19]
    .io_x1(m_114_io_x1),
    .io_x2(m_114_io_x2),
    .io_x3(m_114_io_x3),
    .io_s(m_114_io_s),
    .io_cout(m_114_io_cout)
  );
  Adder m_115 ( // @[MUL.scala 102:19]
    .io_x1(m_115_io_x1),
    .io_x2(m_115_io_x2),
    .io_x3(m_115_io_x3),
    .io_s(m_115_io_s),
    .io_cout(m_115_io_cout)
  );
  Adder m_116 ( // @[MUL.scala 102:19]
    .io_x1(m_116_io_x1),
    .io_x2(m_116_io_x2),
    .io_x3(m_116_io_x3),
    .io_s(m_116_io_s),
    .io_cout(m_116_io_cout)
  );
  Adder m_117 ( // @[MUL.scala 102:19]
    .io_x1(m_117_io_x1),
    .io_x2(m_117_io_x2),
    .io_x3(m_117_io_x3),
    .io_s(m_117_io_s),
    .io_cout(m_117_io_cout)
  );
  Adder m_118 ( // @[MUL.scala 102:19]
    .io_x1(m_118_io_x1),
    .io_x2(m_118_io_x2),
    .io_x3(m_118_io_x3),
    .io_s(m_118_io_s),
    .io_cout(m_118_io_cout)
  );
  Adder m_119 ( // @[MUL.scala 102:19]
    .io_x1(m_119_io_x1),
    .io_x2(m_119_io_x2),
    .io_x3(m_119_io_x3),
    .io_s(m_119_io_s),
    .io_cout(m_119_io_cout)
  );
  Adder m_120 ( // @[MUL.scala 102:19]
    .io_x1(m_120_io_x1),
    .io_x2(m_120_io_x2),
    .io_x3(m_120_io_x3),
    .io_s(m_120_io_s),
    .io_cout(m_120_io_cout)
  );
  Adder m_121 ( // @[MUL.scala 102:19]
    .io_x1(m_121_io_x1),
    .io_x2(m_121_io_x2),
    .io_x3(m_121_io_x3),
    .io_s(m_121_io_s),
    .io_cout(m_121_io_cout)
  );
  Adder m_122 ( // @[MUL.scala 102:19]
    .io_x1(m_122_io_x1),
    .io_x2(m_122_io_x2),
    .io_x3(m_122_io_x3),
    .io_s(m_122_io_s),
    .io_cout(m_122_io_cout)
  );
  Adder m_123 ( // @[MUL.scala 102:19]
    .io_x1(m_123_io_x1),
    .io_x2(m_123_io_x2),
    .io_x3(m_123_io_x3),
    .io_s(m_123_io_s),
    .io_cout(m_123_io_cout)
  );
  Adder m_124 ( // @[MUL.scala 102:19]
    .io_x1(m_124_io_x1),
    .io_x2(m_124_io_x2),
    .io_x3(m_124_io_x3),
    .io_s(m_124_io_s),
    .io_cout(m_124_io_cout)
  );
  Adder m_125 ( // @[MUL.scala 102:19]
    .io_x1(m_125_io_x1),
    .io_x2(m_125_io_x2),
    .io_x3(m_125_io_x3),
    .io_s(m_125_io_s),
    .io_cout(m_125_io_cout)
  );
  Adder m_126 ( // @[MUL.scala 102:19]
    .io_x1(m_126_io_x1),
    .io_x2(m_126_io_x2),
    .io_x3(m_126_io_x3),
    .io_s(m_126_io_s),
    .io_cout(m_126_io_cout)
  );
  Adder m_127 ( // @[MUL.scala 102:19]
    .io_x1(m_127_io_x1),
    .io_x2(m_127_io_x2),
    .io_x3(m_127_io_x3),
    .io_s(m_127_io_s),
    .io_cout(m_127_io_cout)
  );
  Half_Adder m_128 ( // @[MUL.scala 124:19]
    .io_in_0(m_128_io_in_0),
    .io_in_1(m_128_io_in_1),
    .io_out_0(m_128_io_out_0),
    .io_out_1(m_128_io_out_1)
  );
  Adder m_129 ( // @[MUL.scala 102:19]
    .io_x1(m_129_io_x1),
    .io_x2(m_129_io_x2),
    .io_x3(m_129_io_x3),
    .io_s(m_129_io_s),
    .io_cout(m_129_io_cout)
  );
  Adder m_130 ( // @[MUL.scala 102:19]
    .io_x1(m_130_io_x1),
    .io_x2(m_130_io_x2),
    .io_x3(m_130_io_x3),
    .io_s(m_130_io_s),
    .io_cout(m_130_io_cout)
  );
  Adder m_131 ( // @[MUL.scala 102:19]
    .io_x1(m_131_io_x1),
    .io_x2(m_131_io_x2),
    .io_x3(m_131_io_x3),
    .io_s(m_131_io_s),
    .io_cout(m_131_io_cout)
  );
  Adder m_132 ( // @[MUL.scala 102:19]
    .io_x1(m_132_io_x1),
    .io_x2(m_132_io_x2),
    .io_x3(m_132_io_x3),
    .io_s(m_132_io_s),
    .io_cout(m_132_io_cout)
  );
  Adder m_133 ( // @[MUL.scala 102:19]
    .io_x1(m_133_io_x1),
    .io_x2(m_133_io_x2),
    .io_x3(m_133_io_x3),
    .io_s(m_133_io_s),
    .io_cout(m_133_io_cout)
  );
  Half_Adder m_134 ( // @[MUL.scala 124:19]
    .io_in_0(m_134_io_in_0),
    .io_in_1(m_134_io_in_1),
    .io_out_0(m_134_io_out_0),
    .io_out_1(m_134_io_out_1)
  );
  Adder m_135 ( // @[MUL.scala 102:19]
    .io_x1(m_135_io_x1),
    .io_x2(m_135_io_x2),
    .io_x3(m_135_io_x3),
    .io_s(m_135_io_s),
    .io_cout(m_135_io_cout)
  );
  Adder m_136 ( // @[MUL.scala 102:19]
    .io_x1(m_136_io_x1),
    .io_x2(m_136_io_x2),
    .io_x3(m_136_io_x3),
    .io_s(m_136_io_s),
    .io_cout(m_136_io_cout)
  );
  Adder m_137 ( // @[MUL.scala 102:19]
    .io_x1(m_137_io_x1),
    .io_x2(m_137_io_x2),
    .io_x3(m_137_io_x3),
    .io_s(m_137_io_s),
    .io_cout(m_137_io_cout)
  );
  Adder m_138 ( // @[MUL.scala 102:19]
    .io_x1(m_138_io_x1),
    .io_x2(m_138_io_x2),
    .io_x3(m_138_io_x3),
    .io_s(m_138_io_s),
    .io_cout(m_138_io_cout)
  );
  Adder m_139 ( // @[MUL.scala 102:19]
    .io_x1(m_139_io_x1),
    .io_x2(m_139_io_x2),
    .io_x3(m_139_io_x3),
    .io_s(m_139_io_s),
    .io_cout(m_139_io_cout)
  );
  Adder m_140 ( // @[MUL.scala 102:19]
    .io_x1(m_140_io_x1),
    .io_x2(m_140_io_x2),
    .io_x3(m_140_io_x3),
    .io_s(m_140_io_s),
    .io_cout(m_140_io_cout)
  );
  Adder m_141 ( // @[MUL.scala 102:19]
    .io_x1(m_141_io_x1),
    .io_x2(m_141_io_x2),
    .io_x3(m_141_io_x3),
    .io_s(m_141_io_s),
    .io_cout(m_141_io_cout)
  );
  Adder m_142 ( // @[MUL.scala 102:19]
    .io_x1(m_142_io_x1),
    .io_x2(m_142_io_x2),
    .io_x3(m_142_io_x3),
    .io_s(m_142_io_s),
    .io_cout(m_142_io_cout)
  );
  Adder m_143 ( // @[MUL.scala 102:19]
    .io_x1(m_143_io_x1),
    .io_x2(m_143_io_x2),
    .io_x3(m_143_io_x3),
    .io_s(m_143_io_s),
    .io_cout(m_143_io_cout)
  );
  Adder m_144 ( // @[MUL.scala 102:19]
    .io_x1(m_144_io_x1),
    .io_x2(m_144_io_x2),
    .io_x3(m_144_io_x3),
    .io_s(m_144_io_s),
    .io_cout(m_144_io_cout)
  );
  Adder m_145 ( // @[MUL.scala 102:19]
    .io_x1(m_145_io_x1),
    .io_x2(m_145_io_x2),
    .io_x3(m_145_io_x3),
    .io_s(m_145_io_s),
    .io_cout(m_145_io_cout)
  );
  Adder m_146 ( // @[MUL.scala 102:19]
    .io_x1(m_146_io_x1),
    .io_x2(m_146_io_x2),
    .io_x3(m_146_io_x3),
    .io_s(m_146_io_s),
    .io_cout(m_146_io_cout)
  );
  Adder m_147 ( // @[MUL.scala 102:19]
    .io_x1(m_147_io_x1),
    .io_x2(m_147_io_x2),
    .io_x3(m_147_io_x3),
    .io_s(m_147_io_s),
    .io_cout(m_147_io_cout)
  );
  Adder m_148 ( // @[MUL.scala 102:19]
    .io_x1(m_148_io_x1),
    .io_x2(m_148_io_x2),
    .io_x3(m_148_io_x3),
    .io_s(m_148_io_s),
    .io_cout(m_148_io_cout)
  );
  Adder m_149 ( // @[MUL.scala 102:19]
    .io_x1(m_149_io_x1),
    .io_x2(m_149_io_x2),
    .io_x3(m_149_io_x3),
    .io_s(m_149_io_s),
    .io_cout(m_149_io_cout)
  );
  Adder m_150 ( // @[MUL.scala 102:19]
    .io_x1(m_150_io_x1),
    .io_x2(m_150_io_x2),
    .io_x3(m_150_io_x3),
    .io_s(m_150_io_s),
    .io_cout(m_150_io_cout)
  );
  Adder m_151 ( // @[MUL.scala 102:19]
    .io_x1(m_151_io_x1),
    .io_x2(m_151_io_x2),
    .io_x3(m_151_io_x3),
    .io_s(m_151_io_s),
    .io_cout(m_151_io_cout)
  );
  Adder m_152 ( // @[MUL.scala 102:19]
    .io_x1(m_152_io_x1),
    .io_x2(m_152_io_x2),
    .io_x3(m_152_io_x3),
    .io_s(m_152_io_s),
    .io_cout(m_152_io_cout)
  );
  Adder m_153 ( // @[MUL.scala 102:19]
    .io_x1(m_153_io_x1),
    .io_x2(m_153_io_x2),
    .io_x3(m_153_io_x3),
    .io_s(m_153_io_s),
    .io_cout(m_153_io_cout)
  );
  Adder m_154 ( // @[MUL.scala 102:19]
    .io_x1(m_154_io_x1),
    .io_x2(m_154_io_x2),
    .io_x3(m_154_io_x3),
    .io_s(m_154_io_s),
    .io_cout(m_154_io_cout)
  );
  Adder m_155 ( // @[MUL.scala 102:19]
    .io_x1(m_155_io_x1),
    .io_x2(m_155_io_x2),
    .io_x3(m_155_io_x3),
    .io_s(m_155_io_s),
    .io_cout(m_155_io_cout)
  );
  Adder m_156 ( // @[MUL.scala 102:19]
    .io_x1(m_156_io_x1),
    .io_x2(m_156_io_x2),
    .io_x3(m_156_io_x3),
    .io_s(m_156_io_s),
    .io_cout(m_156_io_cout)
  );
  Adder m_157 ( // @[MUL.scala 102:19]
    .io_x1(m_157_io_x1),
    .io_x2(m_157_io_x2),
    .io_x3(m_157_io_x3),
    .io_s(m_157_io_s),
    .io_cout(m_157_io_cout)
  );
  Adder m_158 ( // @[MUL.scala 102:19]
    .io_x1(m_158_io_x1),
    .io_x2(m_158_io_x2),
    .io_x3(m_158_io_x3),
    .io_s(m_158_io_s),
    .io_cout(m_158_io_cout)
  );
  Adder m_159 ( // @[MUL.scala 102:19]
    .io_x1(m_159_io_x1),
    .io_x2(m_159_io_x2),
    .io_x3(m_159_io_x3),
    .io_s(m_159_io_s),
    .io_cout(m_159_io_cout)
  );
  Adder m_160 ( // @[MUL.scala 102:19]
    .io_x1(m_160_io_x1),
    .io_x2(m_160_io_x2),
    .io_x3(m_160_io_x3),
    .io_s(m_160_io_s),
    .io_cout(m_160_io_cout)
  );
  Adder m_161 ( // @[MUL.scala 102:19]
    .io_x1(m_161_io_x1),
    .io_x2(m_161_io_x2),
    .io_x3(m_161_io_x3),
    .io_s(m_161_io_s),
    .io_cout(m_161_io_cout)
  );
  Adder m_162 ( // @[MUL.scala 102:19]
    .io_x1(m_162_io_x1),
    .io_x2(m_162_io_x2),
    .io_x3(m_162_io_x3),
    .io_s(m_162_io_s),
    .io_cout(m_162_io_cout)
  );
  Adder m_163 ( // @[MUL.scala 102:19]
    .io_x1(m_163_io_x1),
    .io_x2(m_163_io_x2),
    .io_x3(m_163_io_x3),
    .io_s(m_163_io_s),
    .io_cout(m_163_io_cout)
  );
  Adder m_164 ( // @[MUL.scala 102:19]
    .io_x1(m_164_io_x1),
    .io_x2(m_164_io_x2),
    .io_x3(m_164_io_x3),
    .io_s(m_164_io_s),
    .io_cout(m_164_io_cout)
  );
  Half_Adder m_165 ( // @[MUL.scala 124:19]
    .io_in_0(m_165_io_in_0),
    .io_in_1(m_165_io_in_1),
    .io_out_0(m_165_io_out_0),
    .io_out_1(m_165_io_out_1)
  );
  Adder m_166 ( // @[MUL.scala 102:19]
    .io_x1(m_166_io_x1),
    .io_x2(m_166_io_x2),
    .io_x3(m_166_io_x3),
    .io_s(m_166_io_s),
    .io_cout(m_166_io_cout)
  );
  Adder m_167 ( // @[MUL.scala 102:19]
    .io_x1(m_167_io_x1),
    .io_x2(m_167_io_x2),
    .io_x3(m_167_io_x3),
    .io_s(m_167_io_s),
    .io_cout(m_167_io_cout)
  );
  Adder m_168 ( // @[MUL.scala 102:19]
    .io_x1(m_168_io_x1),
    .io_x2(m_168_io_x2),
    .io_x3(m_168_io_x3),
    .io_s(m_168_io_s),
    .io_cout(m_168_io_cout)
  );
  Adder m_169 ( // @[MUL.scala 102:19]
    .io_x1(m_169_io_x1),
    .io_x2(m_169_io_x2),
    .io_x3(m_169_io_x3),
    .io_s(m_169_io_s),
    .io_cout(m_169_io_cout)
  );
  Adder m_170 ( // @[MUL.scala 102:19]
    .io_x1(m_170_io_x1),
    .io_x2(m_170_io_x2),
    .io_x3(m_170_io_x3),
    .io_s(m_170_io_s),
    .io_cout(m_170_io_cout)
  );
  Adder m_171 ( // @[MUL.scala 102:19]
    .io_x1(m_171_io_x1),
    .io_x2(m_171_io_x2),
    .io_x3(m_171_io_x3),
    .io_s(m_171_io_s),
    .io_cout(m_171_io_cout)
  );
  Half_Adder m_172 ( // @[MUL.scala 124:19]
    .io_in_0(m_172_io_in_0),
    .io_in_1(m_172_io_in_1),
    .io_out_0(m_172_io_out_0),
    .io_out_1(m_172_io_out_1)
  );
  Adder m_173 ( // @[MUL.scala 102:19]
    .io_x1(m_173_io_x1),
    .io_x2(m_173_io_x2),
    .io_x3(m_173_io_x3),
    .io_s(m_173_io_s),
    .io_cout(m_173_io_cout)
  );
  Adder m_174 ( // @[MUL.scala 102:19]
    .io_x1(m_174_io_x1),
    .io_x2(m_174_io_x2),
    .io_x3(m_174_io_x3),
    .io_s(m_174_io_s),
    .io_cout(m_174_io_cout)
  );
  Adder m_175 ( // @[MUL.scala 102:19]
    .io_x1(m_175_io_x1),
    .io_x2(m_175_io_x2),
    .io_x3(m_175_io_x3),
    .io_s(m_175_io_s),
    .io_cout(m_175_io_cout)
  );
  Adder m_176 ( // @[MUL.scala 102:19]
    .io_x1(m_176_io_x1),
    .io_x2(m_176_io_x2),
    .io_x3(m_176_io_x3),
    .io_s(m_176_io_s),
    .io_cout(m_176_io_cout)
  );
  Adder m_177 ( // @[MUL.scala 102:19]
    .io_x1(m_177_io_x1),
    .io_x2(m_177_io_x2),
    .io_x3(m_177_io_x3),
    .io_s(m_177_io_s),
    .io_cout(m_177_io_cout)
  );
  Adder m_178 ( // @[MUL.scala 102:19]
    .io_x1(m_178_io_x1),
    .io_x2(m_178_io_x2),
    .io_x3(m_178_io_x3),
    .io_s(m_178_io_s),
    .io_cout(m_178_io_cout)
  );
  Adder m_179 ( // @[MUL.scala 102:19]
    .io_x1(m_179_io_x1),
    .io_x2(m_179_io_x2),
    .io_x3(m_179_io_x3),
    .io_s(m_179_io_s),
    .io_cout(m_179_io_cout)
  );
  Adder m_180 ( // @[MUL.scala 102:19]
    .io_x1(m_180_io_x1),
    .io_x2(m_180_io_x2),
    .io_x3(m_180_io_x3),
    .io_s(m_180_io_s),
    .io_cout(m_180_io_cout)
  );
  Adder m_181 ( // @[MUL.scala 102:19]
    .io_x1(m_181_io_x1),
    .io_x2(m_181_io_x2),
    .io_x3(m_181_io_x3),
    .io_s(m_181_io_s),
    .io_cout(m_181_io_cout)
  );
  Adder m_182 ( // @[MUL.scala 102:19]
    .io_x1(m_182_io_x1),
    .io_x2(m_182_io_x2),
    .io_x3(m_182_io_x3),
    .io_s(m_182_io_s),
    .io_cout(m_182_io_cout)
  );
  Adder m_183 ( // @[MUL.scala 102:19]
    .io_x1(m_183_io_x1),
    .io_x2(m_183_io_x2),
    .io_x3(m_183_io_x3),
    .io_s(m_183_io_s),
    .io_cout(m_183_io_cout)
  );
  Adder m_184 ( // @[MUL.scala 102:19]
    .io_x1(m_184_io_x1),
    .io_x2(m_184_io_x2),
    .io_x3(m_184_io_x3),
    .io_s(m_184_io_s),
    .io_cout(m_184_io_cout)
  );
  Adder m_185 ( // @[MUL.scala 102:19]
    .io_x1(m_185_io_x1),
    .io_x2(m_185_io_x2),
    .io_x3(m_185_io_x3),
    .io_s(m_185_io_s),
    .io_cout(m_185_io_cout)
  );
  Adder m_186 ( // @[MUL.scala 102:19]
    .io_x1(m_186_io_x1),
    .io_x2(m_186_io_x2),
    .io_x3(m_186_io_x3),
    .io_s(m_186_io_s),
    .io_cout(m_186_io_cout)
  );
  Adder m_187 ( // @[MUL.scala 102:19]
    .io_x1(m_187_io_x1),
    .io_x2(m_187_io_x2),
    .io_x3(m_187_io_x3),
    .io_s(m_187_io_s),
    .io_cout(m_187_io_cout)
  );
  Adder m_188 ( // @[MUL.scala 102:19]
    .io_x1(m_188_io_x1),
    .io_x2(m_188_io_x2),
    .io_x3(m_188_io_x3),
    .io_s(m_188_io_s),
    .io_cout(m_188_io_cout)
  );
  Adder m_189 ( // @[MUL.scala 102:19]
    .io_x1(m_189_io_x1),
    .io_x2(m_189_io_x2),
    .io_x3(m_189_io_x3),
    .io_s(m_189_io_s),
    .io_cout(m_189_io_cout)
  );
  Adder m_190 ( // @[MUL.scala 102:19]
    .io_x1(m_190_io_x1),
    .io_x2(m_190_io_x2),
    .io_x3(m_190_io_x3),
    .io_s(m_190_io_s),
    .io_cout(m_190_io_cout)
  );
  Adder m_191 ( // @[MUL.scala 102:19]
    .io_x1(m_191_io_x1),
    .io_x2(m_191_io_x2),
    .io_x3(m_191_io_x3),
    .io_s(m_191_io_s),
    .io_cout(m_191_io_cout)
  );
  Adder m_192 ( // @[MUL.scala 102:19]
    .io_x1(m_192_io_x1),
    .io_x2(m_192_io_x2),
    .io_x3(m_192_io_x3),
    .io_s(m_192_io_s),
    .io_cout(m_192_io_cout)
  );
  Adder m_193 ( // @[MUL.scala 102:19]
    .io_x1(m_193_io_x1),
    .io_x2(m_193_io_x2),
    .io_x3(m_193_io_x3),
    .io_s(m_193_io_s),
    .io_cout(m_193_io_cout)
  );
  Adder m_194 ( // @[MUL.scala 102:19]
    .io_x1(m_194_io_x1),
    .io_x2(m_194_io_x2),
    .io_x3(m_194_io_x3),
    .io_s(m_194_io_s),
    .io_cout(m_194_io_cout)
  );
  Adder m_195 ( // @[MUL.scala 102:19]
    .io_x1(m_195_io_x1),
    .io_x2(m_195_io_x2),
    .io_x3(m_195_io_x3),
    .io_s(m_195_io_s),
    .io_cout(m_195_io_cout)
  );
  Adder m_196 ( // @[MUL.scala 102:19]
    .io_x1(m_196_io_x1),
    .io_x2(m_196_io_x2),
    .io_x3(m_196_io_x3),
    .io_s(m_196_io_s),
    .io_cout(m_196_io_cout)
  );
  Adder m_197 ( // @[MUL.scala 102:19]
    .io_x1(m_197_io_x1),
    .io_x2(m_197_io_x2),
    .io_x3(m_197_io_x3),
    .io_s(m_197_io_s),
    .io_cout(m_197_io_cout)
  );
  Adder m_198 ( // @[MUL.scala 102:19]
    .io_x1(m_198_io_x1),
    .io_x2(m_198_io_x2),
    .io_x3(m_198_io_x3),
    .io_s(m_198_io_s),
    .io_cout(m_198_io_cout)
  );
  Adder m_199 ( // @[MUL.scala 102:19]
    .io_x1(m_199_io_x1),
    .io_x2(m_199_io_x2),
    .io_x3(m_199_io_x3),
    .io_s(m_199_io_s),
    .io_cout(m_199_io_cout)
  );
  Adder m_200 ( // @[MUL.scala 102:19]
    .io_x1(m_200_io_x1),
    .io_x2(m_200_io_x2),
    .io_x3(m_200_io_x3),
    .io_s(m_200_io_s),
    .io_cout(m_200_io_cout)
  );
  Adder m_201 ( // @[MUL.scala 102:19]
    .io_x1(m_201_io_x1),
    .io_x2(m_201_io_x2),
    .io_x3(m_201_io_x3),
    .io_s(m_201_io_s),
    .io_cout(m_201_io_cout)
  );
  Adder m_202 ( // @[MUL.scala 102:19]
    .io_x1(m_202_io_x1),
    .io_x2(m_202_io_x2),
    .io_x3(m_202_io_x3),
    .io_s(m_202_io_s),
    .io_cout(m_202_io_cout)
  );
  Adder m_203 ( // @[MUL.scala 102:19]
    .io_x1(m_203_io_x1),
    .io_x2(m_203_io_x2),
    .io_x3(m_203_io_x3),
    .io_s(m_203_io_s),
    .io_cout(m_203_io_cout)
  );
  Adder m_204 ( // @[MUL.scala 102:19]
    .io_x1(m_204_io_x1),
    .io_x2(m_204_io_x2),
    .io_x3(m_204_io_x3),
    .io_s(m_204_io_s),
    .io_cout(m_204_io_cout)
  );
  Adder m_205 ( // @[MUL.scala 102:19]
    .io_x1(m_205_io_x1),
    .io_x2(m_205_io_x2),
    .io_x3(m_205_io_x3),
    .io_s(m_205_io_s),
    .io_cout(m_205_io_cout)
  );
  Adder m_206 ( // @[MUL.scala 102:19]
    .io_x1(m_206_io_x1),
    .io_x2(m_206_io_x2),
    .io_x3(m_206_io_x3),
    .io_s(m_206_io_s),
    .io_cout(m_206_io_cout)
  );
  Adder m_207 ( // @[MUL.scala 102:19]
    .io_x1(m_207_io_x1),
    .io_x2(m_207_io_x2),
    .io_x3(m_207_io_x3),
    .io_s(m_207_io_s),
    .io_cout(m_207_io_cout)
  );
  Half_Adder m_208 ( // @[MUL.scala 124:19]
    .io_in_0(m_208_io_in_0),
    .io_in_1(m_208_io_in_1),
    .io_out_0(m_208_io_out_0),
    .io_out_1(m_208_io_out_1)
  );
  Adder m_209 ( // @[MUL.scala 102:19]
    .io_x1(m_209_io_x1),
    .io_x2(m_209_io_x2),
    .io_x3(m_209_io_x3),
    .io_s(m_209_io_s),
    .io_cout(m_209_io_cout)
  );
  Adder m_210 ( // @[MUL.scala 102:19]
    .io_x1(m_210_io_x1),
    .io_x2(m_210_io_x2),
    .io_x3(m_210_io_x3),
    .io_s(m_210_io_s),
    .io_cout(m_210_io_cout)
  );
  Adder m_211 ( // @[MUL.scala 102:19]
    .io_x1(m_211_io_x1),
    .io_x2(m_211_io_x2),
    .io_x3(m_211_io_x3),
    .io_s(m_211_io_s),
    .io_cout(m_211_io_cout)
  );
  Adder m_212 ( // @[MUL.scala 102:19]
    .io_x1(m_212_io_x1),
    .io_x2(m_212_io_x2),
    .io_x3(m_212_io_x3),
    .io_s(m_212_io_s),
    .io_cout(m_212_io_cout)
  );
  Adder m_213 ( // @[MUL.scala 102:19]
    .io_x1(m_213_io_x1),
    .io_x2(m_213_io_x2),
    .io_x3(m_213_io_x3),
    .io_s(m_213_io_s),
    .io_cout(m_213_io_cout)
  );
  Adder m_214 ( // @[MUL.scala 102:19]
    .io_x1(m_214_io_x1),
    .io_x2(m_214_io_x2),
    .io_x3(m_214_io_x3),
    .io_s(m_214_io_s),
    .io_cout(m_214_io_cout)
  );
  Adder m_215 ( // @[MUL.scala 102:19]
    .io_x1(m_215_io_x1),
    .io_x2(m_215_io_x2),
    .io_x3(m_215_io_x3),
    .io_s(m_215_io_s),
    .io_cout(m_215_io_cout)
  );
  Half_Adder m_216 ( // @[MUL.scala 124:19]
    .io_in_0(m_216_io_in_0),
    .io_in_1(m_216_io_in_1),
    .io_out_0(m_216_io_out_0),
    .io_out_1(m_216_io_out_1)
  );
  Adder m_217 ( // @[MUL.scala 102:19]
    .io_x1(m_217_io_x1),
    .io_x2(m_217_io_x2),
    .io_x3(m_217_io_x3),
    .io_s(m_217_io_s),
    .io_cout(m_217_io_cout)
  );
  Adder m_218 ( // @[MUL.scala 102:19]
    .io_x1(m_218_io_x1),
    .io_x2(m_218_io_x2),
    .io_x3(m_218_io_x3),
    .io_s(m_218_io_s),
    .io_cout(m_218_io_cout)
  );
  Adder m_219 ( // @[MUL.scala 102:19]
    .io_x1(m_219_io_x1),
    .io_x2(m_219_io_x2),
    .io_x3(m_219_io_x3),
    .io_s(m_219_io_s),
    .io_cout(m_219_io_cout)
  );
  Adder m_220 ( // @[MUL.scala 102:19]
    .io_x1(m_220_io_x1),
    .io_x2(m_220_io_x2),
    .io_x3(m_220_io_x3),
    .io_s(m_220_io_s),
    .io_cout(m_220_io_cout)
  );
  Adder m_221 ( // @[MUL.scala 102:19]
    .io_x1(m_221_io_x1),
    .io_x2(m_221_io_x2),
    .io_x3(m_221_io_x3),
    .io_s(m_221_io_s),
    .io_cout(m_221_io_cout)
  );
  Adder m_222 ( // @[MUL.scala 102:19]
    .io_x1(m_222_io_x1),
    .io_x2(m_222_io_x2),
    .io_x3(m_222_io_x3),
    .io_s(m_222_io_s),
    .io_cout(m_222_io_cout)
  );
  Adder m_223 ( // @[MUL.scala 102:19]
    .io_x1(m_223_io_x1),
    .io_x2(m_223_io_x2),
    .io_x3(m_223_io_x3),
    .io_s(m_223_io_s),
    .io_cout(m_223_io_cout)
  );
  Adder m_224 ( // @[MUL.scala 102:19]
    .io_x1(m_224_io_x1),
    .io_x2(m_224_io_x2),
    .io_x3(m_224_io_x3),
    .io_s(m_224_io_s),
    .io_cout(m_224_io_cout)
  );
  Adder m_225 ( // @[MUL.scala 102:19]
    .io_x1(m_225_io_x1),
    .io_x2(m_225_io_x2),
    .io_x3(m_225_io_x3),
    .io_s(m_225_io_s),
    .io_cout(m_225_io_cout)
  );
  Adder m_226 ( // @[MUL.scala 102:19]
    .io_x1(m_226_io_x1),
    .io_x2(m_226_io_x2),
    .io_x3(m_226_io_x3),
    .io_s(m_226_io_s),
    .io_cout(m_226_io_cout)
  );
  Adder m_227 ( // @[MUL.scala 102:19]
    .io_x1(m_227_io_x1),
    .io_x2(m_227_io_x2),
    .io_x3(m_227_io_x3),
    .io_s(m_227_io_s),
    .io_cout(m_227_io_cout)
  );
  Adder m_228 ( // @[MUL.scala 102:19]
    .io_x1(m_228_io_x1),
    .io_x2(m_228_io_x2),
    .io_x3(m_228_io_x3),
    .io_s(m_228_io_s),
    .io_cout(m_228_io_cout)
  );
  Adder m_229 ( // @[MUL.scala 102:19]
    .io_x1(m_229_io_x1),
    .io_x2(m_229_io_x2),
    .io_x3(m_229_io_x3),
    .io_s(m_229_io_s),
    .io_cout(m_229_io_cout)
  );
  Adder m_230 ( // @[MUL.scala 102:19]
    .io_x1(m_230_io_x1),
    .io_x2(m_230_io_x2),
    .io_x3(m_230_io_x3),
    .io_s(m_230_io_s),
    .io_cout(m_230_io_cout)
  );
  Adder m_231 ( // @[MUL.scala 102:19]
    .io_x1(m_231_io_x1),
    .io_x2(m_231_io_x2),
    .io_x3(m_231_io_x3),
    .io_s(m_231_io_s),
    .io_cout(m_231_io_cout)
  );
  Adder m_232 ( // @[MUL.scala 102:19]
    .io_x1(m_232_io_x1),
    .io_x2(m_232_io_x2),
    .io_x3(m_232_io_x3),
    .io_s(m_232_io_s),
    .io_cout(m_232_io_cout)
  );
  Adder m_233 ( // @[MUL.scala 102:19]
    .io_x1(m_233_io_x1),
    .io_x2(m_233_io_x2),
    .io_x3(m_233_io_x3),
    .io_s(m_233_io_s),
    .io_cout(m_233_io_cout)
  );
  Adder m_234 ( // @[MUL.scala 102:19]
    .io_x1(m_234_io_x1),
    .io_x2(m_234_io_x2),
    .io_x3(m_234_io_x3),
    .io_s(m_234_io_s),
    .io_cout(m_234_io_cout)
  );
  Adder m_235 ( // @[MUL.scala 102:19]
    .io_x1(m_235_io_x1),
    .io_x2(m_235_io_x2),
    .io_x3(m_235_io_x3),
    .io_s(m_235_io_s),
    .io_cout(m_235_io_cout)
  );
  Adder m_236 ( // @[MUL.scala 102:19]
    .io_x1(m_236_io_x1),
    .io_x2(m_236_io_x2),
    .io_x3(m_236_io_x3),
    .io_s(m_236_io_s),
    .io_cout(m_236_io_cout)
  );
  Adder m_237 ( // @[MUL.scala 102:19]
    .io_x1(m_237_io_x1),
    .io_x2(m_237_io_x2),
    .io_x3(m_237_io_x3),
    .io_s(m_237_io_s),
    .io_cout(m_237_io_cout)
  );
  Adder m_238 ( // @[MUL.scala 102:19]
    .io_x1(m_238_io_x1),
    .io_x2(m_238_io_x2),
    .io_x3(m_238_io_x3),
    .io_s(m_238_io_s),
    .io_cout(m_238_io_cout)
  );
  Adder m_239 ( // @[MUL.scala 102:19]
    .io_x1(m_239_io_x1),
    .io_x2(m_239_io_x2),
    .io_x3(m_239_io_x3),
    .io_s(m_239_io_s),
    .io_cout(m_239_io_cout)
  );
  Adder m_240 ( // @[MUL.scala 102:19]
    .io_x1(m_240_io_x1),
    .io_x2(m_240_io_x2),
    .io_x3(m_240_io_x3),
    .io_s(m_240_io_s),
    .io_cout(m_240_io_cout)
  );
  Adder m_241 ( // @[MUL.scala 102:19]
    .io_x1(m_241_io_x1),
    .io_x2(m_241_io_x2),
    .io_x3(m_241_io_x3),
    .io_s(m_241_io_s),
    .io_cout(m_241_io_cout)
  );
  Adder m_242 ( // @[MUL.scala 102:19]
    .io_x1(m_242_io_x1),
    .io_x2(m_242_io_x2),
    .io_x3(m_242_io_x3),
    .io_s(m_242_io_s),
    .io_cout(m_242_io_cout)
  );
  Adder m_243 ( // @[MUL.scala 102:19]
    .io_x1(m_243_io_x1),
    .io_x2(m_243_io_x2),
    .io_x3(m_243_io_x3),
    .io_s(m_243_io_s),
    .io_cout(m_243_io_cout)
  );
  Adder m_244 ( // @[MUL.scala 102:19]
    .io_x1(m_244_io_x1),
    .io_x2(m_244_io_x2),
    .io_x3(m_244_io_x3),
    .io_s(m_244_io_s),
    .io_cout(m_244_io_cout)
  );
  Adder m_245 ( // @[MUL.scala 102:19]
    .io_x1(m_245_io_x1),
    .io_x2(m_245_io_x2),
    .io_x3(m_245_io_x3),
    .io_s(m_245_io_s),
    .io_cout(m_245_io_cout)
  );
  Adder m_246 ( // @[MUL.scala 102:19]
    .io_x1(m_246_io_x1),
    .io_x2(m_246_io_x2),
    .io_x3(m_246_io_x3),
    .io_s(m_246_io_s),
    .io_cout(m_246_io_cout)
  );
  Adder m_247 ( // @[MUL.scala 102:19]
    .io_x1(m_247_io_x1),
    .io_x2(m_247_io_x2),
    .io_x3(m_247_io_x3),
    .io_s(m_247_io_s),
    .io_cout(m_247_io_cout)
  );
  Adder m_248 ( // @[MUL.scala 102:19]
    .io_x1(m_248_io_x1),
    .io_x2(m_248_io_x2),
    .io_x3(m_248_io_x3),
    .io_s(m_248_io_s),
    .io_cout(m_248_io_cout)
  );
  Adder m_249 ( // @[MUL.scala 102:19]
    .io_x1(m_249_io_x1),
    .io_x2(m_249_io_x2),
    .io_x3(m_249_io_x3),
    .io_s(m_249_io_s),
    .io_cout(m_249_io_cout)
  );
  Adder m_250 ( // @[MUL.scala 102:19]
    .io_x1(m_250_io_x1),
    .io_x2(m_250_io_x2),
    .io_x3(m_250_io_x3),
    .io_s(m_250_io_s),
    .io_cout(m_250_io_cout)
  );
  Adder m_251 ( // @[MUL.scala 102:19]
    .io_x1(m_251_io_x1),
    .io_x2(m_251_io_x2),
    .io_x3(m_251_io_x3),
    .io_s(m_251_io_s),
    .io_cout(m_251_io_cout)
  );
  Adder m_252 ( // @[MUL.scala 102:19]
    .io_x1(m_252_io_x1),
    .io_x2(m_252_io_x2),
    .io_x3(m_252_io_x3),
    .io_s(m_252_io_s),
    .io_cout(m_252_io_cout)
  );
  Adder m_253 ( // @[MUL.scala 102:19]
    .io_x1(m_253_io_x1),
    .io_x2(m_253_io_x2),
    .io_x3(m_253_io_x3),
    .io_s(m_253_io_s),
    .io_cout(m_253_io_cout)
  );
  Adder m_254 ( // @[MUL.scala 102:19]
    .io_x1(m_254_io_x1),
    .io_x2(m_254_io_x2),
    .io_x3(m_254_io_x3),
    .io_s(m_254_io_s),
    .io_cout(m_254_io_cout)
  );
  Adder m_255 ( // @[MUL.scala 102:19]
    .io_x1(m_255_io_x1),
    .io_x2(m_255_io_x2),
    .io_x3(m_255_io_x3),
    .io_s(m_255_io_s),
    .io_cout(m_255_io_cout)
  );
  Adder m_256 ( // @[MUL.scala 102:19]
    .io_x1(m_256_io_x1),
    .io_x2(m_256_io_x2),
    .io_x3(m_256_io_x3),
    .io_s(m_256_io_s),
    .io_cout(m_256_io_cout)
  );
  Half_Adder m_257 ( // @[MUL.scala 124:19]
    .io_in_0(m_257_io_in_0),
    .io_in_1(m_257_io_in_1),
    .io_out_0(m_257_io_out_0),
    .io_out_1(m_257_io_out_1)
  );
  Adder m_258 ( // @[MUL.scala 102:19]
    .io_x1(m_258_io_x1),
    .io_x2(m_258_io_x2),
    .io_x3(m_258_io_x3),
    .io_s(m_258_io_s),
    .io_cout(m_258_io_cout)
  );
  Adder m_259 ( // @[MUL.scala 102:19]
    .io_x1(m_259_io_x1),
    .io_x2(m_259_io_x2),
    .io_x3(m_259_io_x3),
    .io_s(m_259_io_s),
    .io_cout(m_259_io_cout)
  );
  Adder m_260 ( // @[MUL.scala 102:19]
    .io_x1(m_260_io_x1),
    .io_x2(m_260_io_x2),
    .io_x3(m_260_io_x3),
    .io_s(m_260_io_s),
    .io_cout(m_260_io_cout)
  );
  Adder m_261 ( // @[MUL.scala 102:19]
    .io_x1(m_261_io_x1),
    .io_x2(m_261_io_x2),
    .io_x3(m_261_io_x3),
    .io_s(m_261_io_s),
    .io_cout(m_261_io_cout)
  );
  Adder m_262 ( // @[MUL.scala 102:19]
    .io_x1(m_262_io_x1),
    .io_x2(m_262_io_x2),
    .io_x3(m_262_io_x3),
    .io_s(m_262_io_s),
    .io_cout(m_262_io_cout)
  );
  Adder m_263 ( // @[MUL.scala 102:19]
    .io_x1(m_263_io_x1),
    .io_x2(m_263_io_x2),
    .io_x3(m_263_io_x3),
    .io_s(m_263_io_s),
    .io_cout(m_263_io_cout)
  );
  Adder m_264 ( // @[MUL.scala 102:19]
    .io_x1(m_264_io_x1),
    .io_x2(m_264_io_x2),
    .io_x3(m_264_io_x3),
    .io_s(m_264_io_s),
    .io_cout(m_264_io_cout)
  );
  Adder m_265 ( // @[MUL.scala 102:19]
    .io_x1(m_265_io_x1),
    .io_x2(m_265_io_x2),
    .io_x3(m_265_io_x3),
    .io_s(m_265_io_s),
    .io_cout(m_265_io_cout)
  );
  Half_Adder m_266 ( // @[MUL.scala 124:19]
    .io_in_0(m_266_io_in_0),
    .io_in_1(m_266_io_in_1),
    .io_out_0(m_266_io_out_0),
    .io_out_1(m_266_io_out_1)
  );
  Adder m_267 ( // @[MUL.scala 102:19]
    .io_x1(m_267_io_x1),
    .io_x2(m_267_io_x2),
    .io_x3(m_267_io_x3),
    .io_s(m_267_io_s),
    .io_cout(m_267_io_cout)
  );
  Adder m_268 ( // @[MUL.scala 102:19]
    .io_x1(m_268_io_x1),
    .io_x2(m_268_io_x2),
    .io_x3(m_268_io_x3),
    .io_s(m_268_io_s),
    .io_cout(m_268_io_cout)
  );
  Adder m_269 ( // @[MUL.scala 102:19]
    .io_x1(m_269_io_x1),
    .io_x2(m_269_io_x2),
    .io_x3(m_269_io_x3),
    .io_s(m_269_io_s),
    .io_cout(m_269_io_cout)
  );
  Adder m_270 ( // @[MUL.scala 102:19]
    .io_x1(m_270_io_x1),
    .io_x2(m_270_io_x2),
    .io_x3(m_270_io_x3),
    .io_s(m_270_io_s),
    .io_cout(m_270_io_cout)
  );
  Adder m_271 ( // @[MUL.scala 102:19]
    .io_x1(m_271_io_x1),
    .io_x2(m_271_io_x2),
    .io_x3(m_271_io_x3),
    .io_s(m_271_io_s),
    .io_cout(m_271_io_cout)
  );
  Adder m_272 ( // @[MUL.scala 102:19]
    .io_x1(m_272_io_x1),
    .io_x2(m_272_io_x2),
    .io_x3(m_272_io_x3),
    .io_s(m_272_io_s),
    .io_cout(m_272_io_cout)
  );
  Adder m_273 ( // @[MUL.scala 102:19]
    .io_x1(m_273_io_x1),
    .io_x2(m_273_io_x2),
    .io_x3(m_273_io_x3),
    .io_s(m_273_io_s),
    .io_cout(m_273_io_cout)
  );
  Adder m_274 ( // @[MUL.scala 102:19]
    .io_x1(m_274_io_x1),
    .io_x2(m_274_io_x2),
    .io_x3(m_274_io_x3),
    .io_s(m_274_io_s),
    .io_cout(m_274_io_cout)
  );
  Adder m_275 ( // @[MUL.scala 102:19]
    .io_x1(m_275_io_x1),
    .io_x2(m_275_io_x2),
    .io_x3(m_275_io_x3),
    .io_s(m_275_io_s),
    .io_cout(m_275_io_cout)
  );
  Adder m_276 ( // @[MUL.scala 102:19]
    .io_x1(m_276_io_x1),
    .io_x2(m_276_io_x2),
    .io_x3(m_276_io_x3),
    .io_s(m_276_io_s),
    .io_cout(m_276_io_cout)
  );
  Adder m_277 ( // @[MUL.scala 102:19]
    .io_x1(m_277_io_x1),
    .io_x2(m_277_io_x2),
    .io_x3(m_277_io_x3),
    .io_s(m_277_io_s),
    .io_cout(m_277_io_cout)
  );
  Adder m_278 ( // @[MUL.scala 102:19]
    .io_x1(m_278_io_x1),
    .io_x2(m_278_io_x2),
    .io_x3(m_278_io_x3),
    .io_s(m_278_io_s),
    .io_cout(m_278_io_cout)
  );
  Adder m_279 ( // @[MUL.scala 102:19]
    .io_x1(m_279_io_x1),
    .io_x2(m_279_io_x2),
    .io_x3(m_279_io_x3),
    .io_s(m_279_io_s),
    .io_cout(m_279_io_cout)
  );
  Adder m_280 ( // @[MUL.scala 102:19]
    .io_x1(m_280_io_x1),
    .io_x2(m_280_io_x2),
    .io_x3(m_280_io_x3),
    .io_s(m_280_io_s),
    .io_cout(m_280_io_cout)
  );
  Adder m_281 ( // @[MUL.scala 102:19]
    .io_x1(m_281_io_x1),
    .io_x2(m_281_io_x2),
    .io_x3(m_281_io_x3),
    .io_s(m_281_io_s),
    .io_cout(m_281_io_cout)
  );
  Adder m_282 ( // @[MUL.scala 102:19]
    .io_x1(m_282_io_x1),
    .io_x2(m_282_io_x2),
    .io_x3(m_282_io_x3),
    .io_s(m_282_io_s),
    .io_cout(m_282_io_cout)
  );
  Adder m_283 ( // @[MUL.scala 102:19]
    .io_x1(m_283_io_x1),
    .io_x2(m_283_io_x2),
    .io_x3(m_283_io_x3),
    .io_s(m_283_io_s),
    .io_cout(m_283_io_cout)
  );
  Adder m_284 ( // @[MUL.scala 102:19]
    .io_x1(m_284_io_x1),
    .io_x2(m_284_io_x2),
    .io_x3(m_284_io_x3),
    .io_s(m_284_io_s),
    .io_cout(m_284_io_cout)
  );
  Adder m_285 ( // @[MUL.scala 102:19]
    .io_x1(m_285_io_x1),
    .io_x2(m_285_io_x2),
    .io_x3(m_285_io_x3),
    .io_s(m_285_io_s),
    .io_cout(m_285_io_cout)
  );
  Adder m_286 ( // @[MUL.scala 102:19]
    .io_x1(m_286_io_x1),
    .io_x2(m_286_io_x2),
    .io_x3(m_286_io_x3),
    .io_s(m_286_io_s),
    .io_cout(m_286_io_cout)
  );
  Adder m_287 ( // @[MUL.scala 102:19]
    .io_x1(m_287_io_x1),
    .io_x2(m_287_io_x2),
    .io_x3(m_287_io_x3),
    .io_s(m_287_io_s),
    .io_cout(m_287_io_cout)
  );
  Adder m_288 ( // @[MUL.scala 102:19]
    .io_x1(m_288_io_x1),
    .io_x2(m_288_io_x2),
    .io_x3(m_288_io_x3),
    .io_s(m_288_io_s),
    .io_cout(m_288_io_cout)
  );
  Adder m_289 ( // @[MUL.scala 102:19]
    .io_x1(m_289_io_x1),
    .io_x2(m_289_io_x2),
    .io_x3(m_289_io_x3),
    .io_s(m_289_io_s),
    .io_cout(m_289_io_cout)
  );
  Adder m_290 ( // @[MUL.scala 102:19]
    .io_x1(m_290_io_x1),
    .io_x2(m_290_io_x2),
    .io_x3(m_290_io_x3),
    .io_s(m_290_io_s),
    .io_cout(m_290_io_cout)
  );
  Adder m_291 ( // @[MUL.scala 102:19]
    .io_x1(m_291_io_x1),
    .io_x2(m_291_io_x2),
    .io_x3(m_291_io_x3),
    .io_s(m_291_io_s),
    .io_cout(m_291_io_cout)
  );
  Adder m_292 ( // @[MUL.scala 102:19]
    .io_x1(m_292_io_x1),
    .io_x2(m_292_io_x2),
    .io_x3(m_292_io_x3),
    .io_s(m_292_io_s),
    .io_cout(m_292_io_cout)
  );
  Adder m_293 ( // @[MUL.scala 102:19]
    .io_x1(m_293_io_x1),
    .io_x2(m_293_io_x2),
    .io_x3(m_293_io_x3),
    .io_s(m_293_io_s),
    .io_cout(m_293_io_cout)
  );
  Adder m_294 ( // @[MUL.scala 102:19]
    .io_x1(m_294_io_x1),
    .io_x2(m_294_io_x2),
    .io_x3(m_294_io_x3),
    .io_s(m_294_io_s),
    .io_cout(m_294_io_cout)
  );
  Adder m_295 ( // @[MUL.scala 102:19]
    .io_x1(m_295_io_x1),
    .io_x2(m_295_io_x2),
    .io_x3(m_295_io_x3),
    .io_s(m_295_io_s),
    .io_cout(m_295_io_cout)
  );
  Adder m_296 ( // @[MUL.scala 102:19]
    .io_x1(m_296_io_x1),
    .io_x2(m_296_io_x2),
    .io_x3(m_296_io_x3),
    .io_s(m_296_io_s),
    .io_cout(m_296_io_cout)
  );
  Adder m_297 ( // @[MUL.scala 102:19]
    .io_x1(m_297_io_x1),
    .io_x2(m_297_io_x2),
    .io_x3(m_297_io_x3),
    .io_s(m_297_io_s),
    .io_cout(m_297_io_cout)
  );
  Adder m_298 ( // @[MUL.scala 102:19]
    .io_x1(m_298_io_x1),
    .io_x2(m_298_io_x2),
    .io_x3(m_298_io_x3),
    .io_s(m_298_io_s),
    .io_cout(m_298_io_cout)
  );
  Adder m_299 ( // @[MUL.scala 102:19]
    .io_x1(m_299_io_x1),
    .io_x2(m_299_io_x2),
    .io_x3(m_299_io_x3),
    .io_s(m_299_io_s),
    .io_cout(m_299_io_cout)
  );
  Adder m_300 ( // @[MUL.scala 102:19]
    .io_x1(m_300_io_x1),
    .io_x2(m_300_io_x2),
    .io_x3(m_300_io_x3),
    .io_s(m_300_io_s),
    .io_cout(m_300_io_cout)
  );
  Adder m_301 ( // @[MUL.scala 102:19]
    .io_x1(m_301_io_x1),
    .io_x2(m_301_io_x2),
    .io_x3(m_301_io_x3),
    .io_s(m_301_io_s),
    .io_cout(m_301_io_cout)
  );
  Adder m_302 ( // @[MUL.scala 102:19]
    .io_x1(m_302_io_x1),
    .io_x2(m_302_io_x2),
    .io_x3(m_302_io_x3),
    .io_s(m_302_io_s),
    .io_cout(m_302_io_cout)
  );
  Adder m_303 ( // @[MUL.scala 102:19]
    .io_x1(m_303_io_x1),
    .io_x2(m_303_io_x2),
    .io_x3(m_303_io_x3),
    .io_s(m_303_io_s),
    .io_cout(m_303_io_cout)
  );
  Adder m_304 ( // @[MUL.scala 102:19]
    .io_x1(m_304_io_x1),
    .io_x2(m_304_io_x2),
    .io_x3(m_304_io_x3),
    .io_s(m_304_io_s),
    .io_cout(m_304_io_cout)
  );
  Adder m_305 ( // @[MUL.scala 102:19]
    .io_x1(m_305_io_x1),
    .io_x2(m_305_io_x2),
    .io_x3(m_305_io_x3),
    .io_s(m_305_io_s),
    .io_cout(m_305_io_cout)
  );
  Adder m_306 ( // @[MUL.scala 102:19]
    .io_x1(m_306_io_x1),
    .io_x2(m_306_io_x2),
    .io_x3(m_306_io_x3),
    .io_s(m_306_io_s),
    .io_cout(m_306_io_cout)
  );
  Adder m_307 ( // @[MUL.scala 102:19]
    .io_x1(m_307_io_x1),
    .io_x2(m_307_io_x2),
    .io_x3(m_307_io_x3),
    .io_s(m_307_io_s),
    .io_cout(m_307_io_cout)
  );
  Adder m_308 ( // @[MUL.scala 102:19]
    .io_x1(m_308_io_x1),
    .io_x2(m_308_io_x2),
    .io_x3(m_308_io_x3),
    .io_s(m_308_io_s),
    .io_cout(m_308_io_cout)
  );
  Adder m_309 ( // @[MUL.scala 102:19]
    .io_x1(m_309_io_x1),
    .io_x2(m_309_io_x2),
    .io_x3(m_309_io_x3),
    .io_s(m_309_io_s),
    .io_cout(m_309_io_cout)
  );
  Adder m_310 ( // @[MUL.scala 102:19]
    .io_x1(m_310_io_x1),
    .io_x2(m_310_io_x2),
    .io_x3(m_310_io_x3),
    .io_s(m_310_io_s),
    .io_cout(m_310_io_cout)
  );
  Adder m_311 ( // @[MUL.scala 102:19]
    .io_x1(m_311_io_x1),
    .io_x2(m_311_io_x2),
    .io_x3(m_311_io_x3),
    .io_s(m_311_io_s),
    .io_cout(m_311_io_cout)
  );
  Half_Adder m_312 ( // @[MUL.scala 124:19]
    .io_in_0(m_312_io_in_0),
    .io_in_1(m_312_io_in_1),
    .io_out_0(m_312_io_out_0),
    .io_out_1(m_312_io_out_1)
  );
  Adder m_313 ( // @[MUL.scala 102:19]
    .io_x1(m_313_io_x1),
    .io_x2(m_313_io_x2),
    .io_x3(m_313_io_x3),
    .io_s(m_313_io_s),
    .io_cout(m_313_io_cout)
  );
  Adder m_314 ( // @[MUL.scala 102:19]
    .io_x1(m_314_io_x1),
    .io_x2(m_314_io_x2),
    .io_x3(m_314_io_x3),
    .io_s(m_314_io_s),
    .io_cout(m_314_io_cout)
  );
  Adder m_315 ( // @[MUL.scala 102:19]
    .io_x1(m_315_io_x1),
    .io_x2(m_315_io_x2),
    .io_x3(m_315_io_x3),
    .io_s(m_315_io_s),
    .io_cout(m_315_io_cout)
  );
  Adder m_316 ( // @[MUL.scala 102:19]
    .io_x1(m_316_io_x1),
    .io_x2(m_316_io_x2),
    .io_x3(m_316_io_x3),
    .io_s(m_316_io_s),
    .io_cout(m_316_io_cout)
  );
  Adder m_317 ( // @[MUL.scala 102:19]
    .io_x1(m_317_io_x1),
    .io_x2(m_317_io_x2),
    .io_x3(m_317_io_x3),
    .io_s(m_317_io_s),
    .io_cout(m_317_io_cout)
  );
  Adder m_318 ( // @[MUL.scala 102:19]
    .io_x1(m_318_io_x1),
    .io_x2(m_318_io_x2),
    .io_x3(m_318_io_x3),
    .io_s(m_318_io_s),
    .io_cout(m_318_io_cout)
  );
  Adder m_319 ( // @[MUL.scala 102:19]
    .io_x1(m_319_io_x1),
    .io_x2(m_319_io_x2),
    .io_x3(m_319_io_x3),
    .io_s(m_319_io_s),
    .io_cout(m_319_io_cout)
  );
  Adder m_320 ( // @[MUL.scala 102:19]
    .io_x1(m_320_io_x1),
    .io_x2(m_320_io_x2),
    .io_x3(m_320_io_x3),
    .io_s(m_320_io_s),
    .io_cout(m_320_io_cout)
  );
  Adder m_321 ( // @[MUL.scala 102:19]
    .io_x1(m_321_io_x1),
    .io_x2(m_321_io_x2),
    .io_x3(m_321_io_x3),
    .io_s(m_321_io_s),
    .io_cout(m_321_io_cout)
  );
  Half_Adder m_322 ( // @[MUL.scala 124:19]
    .io_in_0(m_322_io_in_0),
    .io_in_1(m_322_io_in_1),
    .io_out_0(m_322_io_out_0),
    .io_out_1(m_322_io_out_1)
  );
  Adder m_323 ( // @[MUL.scala 102:19]
    .io_x1(m_323_io_x1),
    .io_x2(m_323_io_x2),
    .io_x3(m_323_io_x3),
    .io_s(m_323_io_s),
    .io_cout(m_323_io_cout)
  );
  Adder m_324 ( // @[MUL.scala 102:19]
    .io_x1(m_324_io_x1),
    .io_x2(m_324_io_x2),
    .io_x3(m_324_io_x3),
    .io_s(m_324_io_s),
    .io_cout(m_324_io_cout)
  );
  Adder m_325 ( // @[MUL.scala 102:19]
    .io_x1(m_325_io_x1),
    .io_x2(m_325_io_x2),
    .io_x3(m_325_io_x3),
    .io_s(m_325_io_s),
    .io_cout(m_325_io_cout)
  );
  Adder m_326 ( // @[MUL.scala 102:19]
    .io_x1(m_326_io_x1),
    .io_x2(m_326_io_x2),
    .io_x3(m_326_io_x3),
    .io_s(m_326_io_s),
    .io_cout(m_326_io_cout)
  );
  Adder m_327 ( // @[MUL.scala 102:19]
    .io_x1(m_327_io_x1),
    .io_x2(m_327_io_x2),
    .io_x3(m_327_io_x3),
    .io_s(m_327_io_s),
    .io_cout(m_327_io_cout)
  );
  Adder m_328 ( // @[MUL.scala 102:19]
    .io_x1(m_328_io_x1),
    .io_x2(m_328_io_x2),
    .io_x3(m_328_io_x3),
    .io_s(m_328_io_s),
    .io_cout(m_328_io_cout)
  );
  Adder m_329 ( // @[MUL.scala 102:19]
    .io_x1(m_329_io_x1),
    .io_x2(m_329_io_x2),
    .io_x3(m_329_io_x3),
    .io_s(m_329_io_s),
    .io_cout(m_329_io_cout)
  );
  Adder m_330 ( // @[MUL.scala 102:19]
    .io_x1(m_330_io_x1),
    .io_x2(m_330_io_x2),
    .io_x3(m_330_io_x3),
    .io_s(m_330_io_s),
    .io_cout(m_330_io_cout)
  );
  Adder m_331 ( // @[MUL.scala 102:19]
    .io_x1(m_331_io_x1),
    .io_x2(m_331_io_x2),
    .io_x3(m_331_io_x3),
    .io_s(m_331_io_s),
    .io_cout(m_331_io_cout)
  );
  Adder m_332 ( // @[MUL.scala 102:19]
    .io_x1(m_332_io_x1),
    .io_x2(m_332_io_x2),
    .io_x3(m_332_io_x3),
    .io_s(m_332_io_s),
    .io_cout(m_332_io_cout)
  );
  Adder m_333 ( // @[MUL.scala 102:19]
    .io_x1(m_333_io_x1),
    .io_x2(m_333_io_x2),
    .io_x3(m_333_io_x3),
    .io_s(m_333_io_s),
    .io_cout(m_333_io_cout)
  );
  Adder m_334 ( // @[MUL.scala 102:19]
    .io_x1(m_334_io_x1),
    .io_x2(m_334_io_x2),
    .io_x3(m_334_io_x3),
    .io_s(m_334_io_s),
    .io_cout(m_334_io_cout)
  );
  Adder m_335 ( // @[MUL.scala 102:19]
    .io_x1(m_335_io_x1),
    .io_x2(m_335_io_x2),
    .io_x3(m_335_io_x3),
    .io_s(m_335_io_s),
    .io_cout(m_335_io_cout)
  );
  Adder m_336 ( // @[MUL.scala 102:19]
    .io_x1(m_336_io_x1),
    .io_x2(m_336_io_x2),
    .io_x3(m_336_io_x3),
    .io_s(m_336_io_s),
    .io_cout(m_336_io_cout)
  );
  Adder m_337 ( // @[MUL.scala 102:19]
    .io_x1(m_337_io_x1),
    .io_x2(m_337_io_x2),
    .io_x3(m_337_io_x3),
    .io_s(m_337_io_s),
    .io_cout(m_337_io_cout)
  );
  Adder m_338 ( // @[MUL.scala 102:19]
    .io_x1(m_338_io_x1),
    .io_x2(m_338_io_x2),
    .io_x3(m_338_io_x3),
    .io_s(m_338_io_s),
    .io_cout(m_338_io_cout)
  );
  Adder m_339 ( // @[MUL.scala 102:19]
    .io_x1(m_339_io_x1),
    .io_x2(m_339_io_x2),
    .io_x3(m_339_io_x3),
    .io_s(m_339_io_s),
    .io_cout(m_339_io_cout)
  );
  Adder m_340 ( // @[MUL.scala 102:19]
    .io_x1(m_340_io_x1),
    .io_x2(m_340_io_x2),
    .io_x3(m_340_io_x3),
    .io_s(m_340_io_s),
    .io_cout(m_340_io_cout)
  );
  Adder m_341 ( // @[MUL.scala 102:19]
    .io_x1(m_341_io_x1),
    .io_x2(m_341_io_x2),
    .io_x3(m_341_io_x3),
    .io_s(m_341_io_s),
    .io_cout(m_341_io_cout)
  );
  Adder m_342 ( // @[MUL.scala 102:19]
    .io_x1(m_342_io_x1),
    .io_x2(m_342_io_x2),
    .io_x3(m_342_io_x3),
    .io_s(m_342_io_s),
    .io_cout(m_342_io_cout)
  );
  Adder m_343 ( // @[MUL.scala 102:19]
    .io_x1(m_343_io_x1),
    .io_x2(m_343_io_x2),
    .io_x3(m_343_io_x3),
    .io_s(m_343_io_s),
    .io_cout(m_343_io_cout)
  );
  Adder m_344 ( // @[MUL.scala 102:19]
    .io_x1(m_344_io_x1),
    .io_x2(m_344_io_x2),
    .io_x3(m_344_io_x3),
    .io_s(m_344_io_s),
    .io_cout(m_344_io_cout)
  );
  Adder m_345 ( // @[MUL.scala 102:19]
    .io_x1(m_345_io_x1),
    .io_x2(m_345_io_x2),
    .io_x3(m_345_io_x3),
    .io_s(m_345_io_s),
    .io_cout(m_345_io_cout)
  );
  Adder m_346 ( // @[MUL.scala 102:19]
    .io_x1(m_346_io_x1),
    .io_x2(m_346_io_x2),
    .io_x3(m_346_io_x3),
    .io_s(m_346_io_s),
    .io_cout(m_346_io_cout)
  );
  Adder m_347 ( // @[MUL.scala 102:19]
    .io_x1(m_347_io_x1),
    .io_x2(m_347_io_x2),
    .io_x3(m_347_io_x3),
    .io_s(m_347_io_s),
    .io_cout(m_347_io_cout)
  );
  Adder m_348 ( // @[MUL.scala 102:19]
    .io_x1(m_348_io_x1),
    .io_x2(m_348_io_x2),
    .io_x3(m_348_io_x3),
    .io_s(m_348_io_s),
    .io_cout(m_348_io_cout)
  );
  Adder m_349 ( // @[MUL.scala 102:19]
    .io_x1(m_349_io_x1),
    .io_x2(m_349_io_x2),
    .io_x3(m_349_io_x3),
    .io_s(m_349_io_s),
    .io_cout(m_349_io_cout)
  );
  Adder m_350 ( // @[MUL.scala 102:19]
    .io_x1(m_350_io_x1),
    .io_x2(m_350_io_x2),
    .io_x3(m_350_io_x3),
    .io_s(m_350_io_s),
    .io_cout(m_350_io_cout)
  );
  Adder m_351 ( // @[MUL.scala 102:19]
    .io_x1(m_351_io_x1),
    .io_x2(m_351_io_x2),
    .io_x3(m_351_io_x3),
    .io_s(m_351_io_s),
    .io_cout(m_351_io_cout)
  );
  Adder m_352 ( // @[MUL.scala 102:19]
    .io_x1(m_352_io_x1),
    .io_x2(m_352_io_x2),
    .io_x3(m_352_io_x3),
    .io_s(m_352_io_s),
    .io_cout(m_352_io_cout)
  );
  Adder m_353 ( // @[MUL.scala 102:19]
    .io_x1(m_353_io_x1),
    .io_x2(m_353_io_x2),
    .io_x3(m_353_io_x3),
    .io_s(m_353_io_s),
    .io_cout(m_353_io_cout)
  );
  Adder m_354 ( // @[MUL.scala 102:19]
    .io_x1(m_354_io_x1),
    .io_x2(m_354_io_x2),
    .io_x3(m_354_io_x3),
    .io_s(m_354_io_s),
    .io_cout(m_354_io_cout)
  );
  Adder m_355 ( // @[MUL.scala 102:19]
    .io_x1(m_355_io_x1),
    .io_x2(m_355_io_x2),
    .io_x3(m_355_io_x3),
    .io_s(m_355_io_s),
    .io_cout(m_355_io_cout)
  );
  Adder m_356 ( // @[MUL.scala 102:19]
    .io_x1(m_356_io_x1),
    .io_x2(m_356_io_x2),
    .io_x3(m_356_io_x3),
    .io_s(m_356_io_s),
    .io_cout(m_356_io_cout)
  );
  Adder m_357 ( // @[MUL.scala 102:19]
    .io_x1(m_357_io_x1),
    .io_x2(m_357_io_x2),
    .io_x3(m_357_io_x3),
    .io_s(m_357_io_s),
    .io_cout(m_357_io_cout)
  );
  Adder m_358 ( // @[MUL.scala 102:19]
    .io_x1(m_358_io_x1),
    .io_x2(m_358_io_x2),
    .io_x3(m_358_io_x3),
    .io_s(m_358_io_s),
    .io_cout(m_358_io_cout)
  );
  Adder m_359 ( // @[MUL.scala 102:19]
    .io_x1(m_359_io_x1),
    .io_x2(m_359_io_x2),
    .io_x3(m_359_io_x3),
    .io_s(m_359_io_s),
    .io_cout(m_359_io_cout)
  );
  Adder m_360 ( // @[MUL.scala 102:19]
    .io_x1(m_360_io_x1),
    .io_x2(m_360_io_x2),
    .io_x3(m_360_io_x3),
    .io_s(m_360_io_s),
    .io_cout(m_360_io_cout)
  );
  Adder m_361 ( // @[MUL.scala 102:19]
    .io_x1(m_361_io_x1),
    .io_x2(m_361_io_x2),
    .io_x3(m_361_io_x3),
    .io_s(m_361_io_s),
    .io_cout(m_361_io_cout)
  );
  Adder m_362 ( // @[MUL.scala 102:19]
    .io_x1(m_362_io_x1),
    .io_x2(m_362_io_x2),
    .io_x3(m_362_io_x3),
    .io_s(m_362_io_s),
    .io_cout(m_362_io_cout)
  );
  Adder m_363 ( // @[MUL.scala 102:19]
    .io_x1(m_363_io_x1),
    .io_x2(m_363_io_x2),
    .io_x3(m_363_io_x3),
    .io_s(m_363_io_s),
    .io_cout(m_363_io_cout)
  );
  Adder m_364 ( // @[MUL.scala 102:19]
    .io_x1(m_364_io_x1),
    .io_x2(m_364_io_x2),
    .io_x3(m_364_io_x3),
    .io_s(m_364_io_s),
    .io_cout(m_364_io_cout)
  );
  Adder m_365 ( // @[MUL.scala 102:19]
    .io_x1(m_365_io_x1),
    .io_x2(m_365_io_x2),
    .io_x3(m_365_io_x3),
    .io_s(m_365_io_s),
    .io_cout(m_365_io_cout)
  );
  Adder m_366 ( // @[MUL.scala 102:19]
    .io_x1(m_366_io_x1),
    .io_x2(m_366_io_x2),
    .io_x3(m_366_io_x3),
    .io_s(m_366_io_s),
    .io_cout(m_366_io_cout)
  );
  Adder m_367 ( // @[MUL.scala 102:19]
    .io_x1(m_367_io_x1),
    .io_x2(m_367_io_x2),
    .io_x3(m_367_io_x3),
    .io_s(m_367_io_s),
    .io_cout(m_367_io_cout)
  );
  Adder m_368 ( // @[MUL.scala 102:19]
    .io_x1(m_368_io_x1),
    .io_x2(m_368_io_x2),
    .io_x3(m_368_io_x3),
    .io_s(m_368_io_s),
    .io_cout(m_368_io_cout)
  );
  Adder m_369 ( // @[MUL.scala 102:19]
    .io_x1(m_369_io_x1),
    .io_x2(m_369_io_x2),
    .io_x3(m_369_io_x3),
    .io_s(m_369_io_s),
    .io_cout(m_369_io_cout)
  );
  Adder m_370 ( // @[MUL.scala 102:19]
    .io_x1(m_370_io_x1),
    .io_x2(m_370_io_x2),
    .io_x3(m_370_io_x3),
    .io_s(m_370_io_s),
    .io_cout(m_370_io_cout)
  );
  Adder m_371 ( // @[MUL.scala 102:19]
    .io_x1(m_371_io_x1),
    .io_x2(m_371_io_x2),
    .io_x3(m_371_io_x3),
    .io_s(m_371_io_s),
    .io_cout(m_371_io_cout)
  );
  Adder m_372 ( // @[MUL.scala 102:19]
    .io_x1(m_372_io_x1),
    .io_x2(m_372_io_x2),
    .io_x3(m_372_io_x3),
    .io_s(m_372_io_s),
    .io_cout(m_372_io_cout)
  );
  Half_Adder m_373 ( // @[MUL.scala 124:19]
    .io_in_0(m_373_io_in_0),
    .io_in_1(m_373_io_in_1),
    .io_out_0(m_373_io_out_0),
    .io_out_1(m_373_io_out_1)
  );
  Adder m_374 ( // @[MUL.scala 102:19]
    .io_x1(m_374_io_x1),
    .io_x2(m_374_io_x2),
    .io_x3(m_374_io_x3),
    .io_s(m_374_io_s),
    .io_cout(m_374_io_cout)
  );
  Adder m_375 ( // @[MUL.scala 102:19]
    .io_x1(m_375_io_x1),
    .io_x2(m_375_io_x2),
    .io_x3(m_375_io_x3),
    .io_s(m_375_io_s),
    .io_cout(m_375_io_cout)
  );
  Adder m_376 ( // @[MUL.scala 102:19]
    .io_x1(m_376_io_x1),
    .io_x2(m_376_io_x2),
    .io_x3(m_376_io_x3),
    .io_s(m_376_io_s),
    .io_cout(m_376_io_cout)
  );
  Adder m_377 ( // @[MUL.scala 102:19]
    .io_x1(m_377_io_x1),
    .io_x2(m_377_io_x2),
    .io_x3(m_377_io_x3),
    .io_s(m_377_io_s),
    .io_cout(m_377_io_cout)
  );
  Adder m_378 ( // @[MUL.scala 102:19]
    .io_x1(m_378_io_x1),
    .io_x2(m_378_io_x2),
    .io_x3(m_378_io_x3),
    .io_s(m_378_io_s),
    .io_cout(m_378_io_cout)
  );
  Adder m_379 ( // @[MUL.scala 102:19]
    .io_x1(m_379_io_x1),
    .io_x2(m_379_io_x2),
    .io_x3(m_379_io_x3),
    .io_s(m_379_io_s),
    .io_cout(m_379_io_cout)
  );
  Adder m_380 ( // @[MUL.scala 102:19]
    .io_x1(m_380_io_x1),
    .io_x2(m_380_io_x2),
    .io_x3(m_380_io_x3),
    .io_s(m_380_io_s),
    .io_cout(m_380_io_cout)
  );
  Adder m_381 ( // @[MUL.scala 102:19]
    .io_x1(m_381_io_x1),
    .io_x2(m_381_io_x2),
    .io_x3(m_381_io_x3),
    .io_s(m_381_io_s),
    .io_cout(m_381_io_cout)
  );
  Adder m_382 ( // @[MUL.scala 102:19]
    .io_x1(m_382_io_x1),
    .io_x2(m_382_io_x2),
    .io_x3(m_382_io_x3),
    .io_s(m_382_io_s),
    .io_cout(m_382_io_cout)
  );
  Adder m_383 ( // @[MUL.scala 102:19]
    .io_x1(m_383_io_x1),
    .io_x2(m_383_io_x2),
    .io_x3(m_383_io_x3),
    .io_s(m_383_io_s),
    .io_cout(m_383_io_cout)
  );
  Half_Adder m_384 ( // @[MUL.scala 124:19]
    .io_in_0(m_384_io_in_0),
    .io_in_1(m_384_io_in_1),
    .io_out_0(m_384_io_out_0),
    .io_out_1(m_384_io_out_1)
  );
  Adder m_385 ( // @[MUL.scala 102:19]
    .io_x1(m_385_io_x1),
    .io_x2(m_385_io_x2),
    .io_x3(m_385_io_x3),
    .io_s(m_385_io_s),
    .io_cout(m_385_io_cout)
  );
  Adder m_386 ( // @[MUL.scala 102:19]
    .io_x1(m_386_io_x1),
    .io_x2(m_386_io_x2),
    .io_x3(m_386_io_x3),
    .io_s(m_386_io_s),
    .io_cout(m_386_io_cout)
  );
  Adder m_387 ( // @[MUL.scala 102:19]
    .io_x1(m_387_io_x1),
    .io_x2(m_387_io_x2),
    .io_x3(m_387_io_x3),
    .io_s(m_387_io_s),
    .io_cout(m_387_io_cout)
  );
  Adder m_388 ( // @[MUL.scala 102:19]
    .io_x1(m_388_io_x1),
    .io_x2(m_388_io_x2),
    .io_x3(m_388_io_x3),
    .io_s(m_388_io_s),
    .io_cout(m_388_io_cout)
  );
  Adder m_389 ( // @[MUL.scala 102:19]
    .io_x1(m_389_io_x1),
    .io_x2(m_389_io_x2),
    .io_x3(m_389_io_x3),
    .io_s(m_389_io_s),
    .io_cout(m_389_io_cout)
  );
  Adder m_390 ( // @[MUL.scala 102:19]
    .io_x1(m_390_io_x1),
    .io_x2(m_390_io_x2),
    .io_x3(m_390_io_x3),
    .io_s(m_390_io_s),
    .io_cout(m_390_io_cout)
  );
  Adder m_391 ( // @[MUL.scala 102:19]
    .io_x1(m_391_io_x1),
    .io_x2(m_391_io_x2),
    .io_x3(m_391_io_x3),
    .io_s(m_391_io_s),
    .io_cout(m_391_io_cout)
  );
  Adder m_392 ( // @[MUL.scala 102:19]
    .io_x1(m_392_io_x1),
    .io_x2(m_392_io_x2),
    .io_x3(m_392_io_x3),
    .io_s(m_392_io_s),
    .io_cout(m_392_io_cout)
  );
  Adder m_393 ( // @[MUL.scala 102:19]
    .io_x1(m_393_io_x1),
    .io_x2(m_393_io_x2),
    .io_x3(m_393_io_x3),
    .io_s(m_393_io_s),
    .io_cout(m_393_io_cout)
  );
  Adder m_394 ( // @[MUL.scala 102:19]
    .io_x1(m_394_io_x1),
    .io_x2(m_394_io_x2),
    .io_x3(m_394_io_x3),
    .io_s(m_394_io_s),
    .io_cout(m_394_io_cout)
  );
  Adder m_395 ( // @[MUL.scala 102:19]
    .io_x1(m_395_io_x1),
    .io_x2(m_395_io_x2),
    .io_x3(m_395_io_x3),
    .io_s(m_395_io_s),
    .io_cout(m_395_io_cout)
  );
  Adder m_396 ( // @[MUL.scala 102:19]
    .io_x1(m_396_io_x1),
    .io_x2(m_396_io_x2),
    .io_x3(m_396_io_x3),
    .io_s(m_396_io_s),
    .io_cout(m_396_io_cout)
  );
  Adder m_397 ( // @[MUL.scala 102:19]
    .io_x1(m_397_io_x1),
    .io_x2(m_397_io_x2),
    .io_x3(m_397_io_x3),
    .io_s(m_397_io_s),
    .io_cout(m_397_io_cout)
  );
  Adder m_398 ( // @[MUL.scala 102:19]
    .io_x1(m_398_io_x1),
    .io_x2(m_398_io_x2),
    .io_x3(m_398_io_x3),
    .io_s(m_398_io_s),
    .io_cout(m_398_io_cout)
  );
  Adder m_399 ( // @[MUL.scala 102:19]
    .io_x1(m_399_io_x1),
    .io_x2(m_399_io_x2),
    .io_x3(m_399_io_x3),
    .io_s(m_399_io_s),
    .io_cout(m_399_io_cout)
  );
  Adder m_400 ( // @[MUL.scala 102:19]
    .io_x1(m_400_io_x1),
    .io_x2(m_400_io_x2),
    .io_x3(m_400_io_x3),
    .io_s(m_400_io_s),
    .io_cout(m_400_io_cout)
  );
  Adder m_401 ( // @[MUL.scala 102:19]
    .io_x1(m_401_io_x1),
    .io_x2(m_401_io_x2),
    .io_x3(m_401_io_x3),
    .io_s(m_401_io_s),
    .io_cout(m_401_io_cout)
  );
  Adder m_402 ( // @[MUL.scala 102:19]
    .io_x1(m_402_io_x1),
    .io_x2(m_402_io_x2),
    .io_x3(m_402_io_x3),
    .io_s(m_402_io_s),
    .io_cout(m_402_io_cout)
  );
  Adder m_403 ( // @[MUL.scala 102:19]
    .io_x1(m_403_io_x1),
    .io_x2(m_403_io_x2),
    .io_x3(m_403_io_x3),
    .io_s(m_403_io_s),
    .io_cout(m_403_io_cout)
  );
  Adder m_404 ( // @[MUL.scala 102:19]
    .io_x1(m_404_io_x1),
    .io_x2(m_404_io_x2),
    .io_x3(m_404_io_x3),
    .io_s(m_404_io_s),
    .io_cout(m_404_io_cout)
  );
  Adder m_405 ( // @[MUL.scala 102:19]
    .io_x1(m_405_io_x1),
    .io_x2(m_405_io_x2),
    .io_x3(m_405_io_x3),
    .io_s(m_405_io_s),
    .io_cout(m_405_io_cout)
  );
  Adder m_406 ( // @[MUL.scala 102:19]
    .io_x1(m_406_io_x1),
    .io_x2(m_406_io_x2),
    .io_x3(m_406_io_x3),
    .io_s(m_406_io_s),
    .io_cout(m_406_io_cout)
  );
  Adder m_407 ( // @[MUL.scala 102:19]
    .io_x1(m_407_io_x1),
    .io_x2(m_407_io_x2),
    .io_x3(m_407_io_x3),
    .io_s(m_407_io_s),
    .io_cout(m_407_io_cout)
  );
  Adder m_408 ( // @[MUL.scala 102:19]
    .io_x1(m_408_io_x1),
    .io_x2(m_408_io_x2),
    .io_x3(m_408_io_x3),
    .io_s(m_408_io_s),
    .io_cout(m_408_io_cout)
  );
  Adder m_409 ( // @[MUL.scala 102:19]
    .io_x1(m_409_io_x1),
    .io_x2(m_409_io_x2),
    .io_x3(m_409_io_x3),
    .io_s(m_409_io_s),
    .io_cout(m_409_io_cout)
  );
  Adder m_410 ( // @[MUL.scala 102:19]
    .io_x1(m_410_io_x1),
    .io_x2(m_410_io_x2),
    .io_x3(m_410_io_x3),
    .io_s(m_410_io_s),
    .io_cout(m_410_io_cout)
  );
  Adder m_411 ( // @[MUL.scala 102:19]
    .io_x1(m_411_io_x1),
    .io_x2(m_411_io_x2),
    .io_x3(m_411_io_x3),
    .io_s(m_411_io_s),
    .io_cout(m_411_io_cout)
  );
  Adder m_412 ( // @[MUL.scala 102:19]
    .io_x1(m_412_io_x1),
    .io_x2(m_412_io_x2),
    .io_x3(m_412_io_x3),
    .io_s(m_412_io_s),
    .io_cout(m_412_io_cout)
  );
  Adder m_413 ( // @[MUL.scala 102:19]
    .io_x1(m_413_io_x1),
    .io_x2(m_413_io_x2),
    .io_x3(m_413_io_x3),
    .io_s(m_413_io_s),
    .io_cout(m_413_io_cout)
  );
  Adder m_414 ( // @[MUL.scala 102:19]
    .io_x1(m_414_io_x1),
    .io_x2(m_414_io_x2),
    .io_x3(m_414_io_x3),
    .io_s(m_414_io_s),
    .io_cout(m_414_io_cout)
  );
  Adder m_415 ( // @[MUL.scala 102:19]
    .io_x1(m_415_io_x1),
    .io_x2(m_415_io_x2),
    .io_x3(m_415_io_x3),
    .io_s(m_415_io_s),
    .io_cout(m_415_io_cout)
  );
  Adder m_416 ( // @[MUL.scala 102:19]
    .io_x1(m_416_io_x1),
    .io_x2(m_416_io_x2),
    .io_x3(m_416_io_x3),
    .io_s(m_416_io_s),
    .io_cout(m_416_io_cout)
  );
  Adder m_417 ( // @[MUL.scala 102:19]
    .io_x1(m_417_io_x1),
    .io_x2(m_417_io_x2),
    .io_x3(m_417_io_x3),
    .io_s(m_417_io_s),
    .io_cout(m_417_io_cout)
  );
  Adder m_418 ( // @[MUL.scala 102:19]
    .io_x1(m_418_io_x1),
    .io_x2(m_418_io_x2),
    .io_x3(m_418_io_x3),
    .io_s(m_418_io_s),
    .io_cout(m_418_io_cout)
  );
  Adder m_419 ( // @[MUL.scala 102:19]
    .io_x1(m_419_io_x1),
    .io_x2(m_419_io_x2),
    .io_x3(m_419_io_x3),
    .io_s(m_419_io_s),
    .io_cout(m_419_io_cout)
  );
  Adder m_420 ( // @[MUL.scala 102:19]
    .io_x1(m_420_io_x1),
    .io_x2(m_420_io_x2),
    .io_x3(m_420_io_x3),
    .io_s(m_420_io_s),
    .io_cout(m_420_io_cout)
  );
  Adder m_421 ( // @[MUL.scala 102:19]
    .io_x1(m_421_io_x1),
    .io_x2(m_421_io_x2),
    .io_x3(m_421_io_x3),
    .io_s(m_421_io_s),
    .io_cout(m_421_io_cout)
  );
  Adder m_422 ( // @[MUL.scala 102:19]
    .io_x1(m_422_io_x1),
    .io_x2(m_422_io_x2),
    .io_x3(m_422_io_x3),
    .io_s(m_422_io_s),
    .io_cout(m_422_io_cout)
  );
  Adder m_423 ( // @[MUL.scala 102:19]
    .io_x1(m_423_io_x1),
    .io_x2(m_423_io_x2),
    .io_x3(m_423_io_x3),
    .io_s(m_423_io_s),
    .io_cout(m_423_io_cout)
  );
  Adder m_424 ( // @[MUL.scala 102:19]
    .io_x1(m_424_io_x1),
    .io_x2(m_424_io_x2),
    .io_x3(m_424_io_x3),
    .io_s(m_424_io_s),
    .io_cout(m_424_io_cout)
  );
  Adder m_425 ( // @[MUL.scala 102:19]
    .io_x1(m_425_io_x1),
    .io_x2(m_425_io_x2),
    .io_x3(m_425_io_x3),
    .io_s(m_425_io_s),
    .io_cout(m_425_io_cout)
  );
  Adder m_426 ( // @[MUL.scala 102:19]
    .io_x1(m_426_io_x1),
    .io_x2(m_426_io_x2),
    .io_x3(m_426_io_x3),
    .io_s(m_426_io_s),
    .io_cout(m_426_io_cout)
  );
  Adder m_427 ( // @[MUL.scala 102:19]
    .io_x1(m_427_io_x1),
    .io_x2(m_427_io_x2),
    .io_x3(m_427_io_x3),
    .io_s(m_427_io_s),
    .io_cout(m_427_io_cout)
  );
  Adder m_428 ( // @[MUL.scala 102:19]
    .io_x1(m_428_io_x1),
    .io_x2(m_428_io_x2),
    .io_x3(m_428_io_x3),
    .io_s(m_428_io_s),
    .io_cout(m_428_io_cout)
  );
  Adder m_429 ( // @[MUL.scala 102:19]
    .io_x1(m_429_io_x1),
    .io_x2(m_429_io_x2),
    .io_x3(m_429_io_x3),
    .io_s(m_429_io_s),
    .io_cout(m_429_io_cout)
  );
  Adder m_430 ( // @[MUL.scala 102:19]
    .io_x1(m_430_io_x1),
    .io_x2(m_430_io_x2),
    .io_x3(m_430_io_x3),
    .io_s(m_430_io_s),
    .io_cout(m_430_io_cout)
  );
  Adder m_431 ( // @[MUL.scala 102:19]
    .io_x1(m_431_io_x1),
    .io_x2(m_431_io_x2),
    .io_x3(m_431_io_x3),
    .io_s(m_431_io_s),
    .io_cout(m_431_io_cout)
  );
  Adder m_432 ( // @[MUL.scala 102:19]
    .io_x1(m_432_io_x1),
    .io_x2(m_432_io_x2),
    .io_x3(m_432_io_x3),
    .io_s(m_432_io_s),
    .io_cout(m_432_io_cout)
  );
  Adder m_433 ( // @[MUL.scala 102:19]
    .io_x1(m_433_io_x1),
    .io_x2(m_433_io_x2),
    .io_x3(m_433_io_x3),
    .io_s(m_433_io_s),
    .io_cout(m_433_io_cout)
  );
  Adder m_434 ( // @[MUL.scala 102:19]
    .io_x1(m_434_io_x1),
    .io_x2(m_434_io_x2),
    .io_x3(m_434_io_x3),
    .io_s(m_434_io_s),
    .io_cout(m_434_io_cout)
  );
  Adder m_435 ( // @[MUL.scala 102:19]
    .io_x1(m_435_io_x1),
    .io_x2(m_435_io_x2),
    .io_x3(m_435_io_x3),
    .io_s(m_435_io_s),
    .io_cout(m_435_io_cout)
  );
  Adder m_436 ( // @[MUL.scala 102:19]
    .io_x1(m_436_io_x1),
    .io_x2(m_436_io_x2),
    .io_x3(m_436_io_x3),
    .io_s(m_436_io_s),
    .io_cout(m_436_io_cout)
  );
  Adder m_437 ( // @[MUL.scala 102:19]
    .io_x1(m_437_io_x1),
    .io_x2(m_437_io_x2),
    .io_x3(m_437_io_x3),
    .io_s(m_437_io_s),
    .io_cout(m_437_io_cout)
  );
  Adder m_438 ( // @[MUL.scala 102:19]
    .io_x1(m_438_io_x1),
    .io_x2(m_438_io_x2),
    .io_x3(m_438_io_x3),
    .io_s(m_438_io_s),
    .io_cout(m_438_io_cout)
  );
  Adder m_439 ( // @[MUL.scala 102:19]
    .io_x1(m_439_io_x1),
    .io_x2(m_439_io_x2),
    .io_x3(m_439_io_x3),
    .io_s(m_439_io_s),
    .io_cout(m_439_io_cout)
  );
  Adder m_440 ( // @[MUL.scala 102:19]
    .io_x1(m_440_io_x1),
    .io_x2(m_440_io_x2),
    .io_x3(m_440_io_x3),
    .io_s(m_440_io_s),
    .io_cout(m_440_io_cout)
  );
  Adder m_441 ( // @[MUL.scala 102:19]
    .io_x1(m_441_io_x1),
    .io_x2(m_441_io_x2),
    .io_x3(m_441_io_x3),
    .io_s(m_441_io_s),
    .io_cout(m_441_io_cout)
  );
  Adder m_442 ( // @[MUL.scala 102:19]
    .io_x1(m_442_io_x1),
    .io_x2(m_442_io_x2),
    .io_x3(m_442_io_x3),
    .io_s(m_442_io_s),
    .io_cout(m_442_io_cout)
  );
  Adder m_443 ( // @[MUL.scala 102:19]
    .io_x1(m_443_io_x1),
    .io_x2(m_443_io_x2),
    .io_x3(m_443_io_x3),
    .io_s(m_443_io_s),
    .io_cout(m_443_io_cout)
  );
  Adder m_444 ( // @[MUL.scala 102:19]
    .io_x1(m_444_io_x1),
    .io_x2(m_444_io_x2),
    .io_x3(m_444_io_x3),
    .io_s(m_444_io_s),
    .io_cout(m_444_io_cout)
  );
  Adder m_445 ( // @[MUL.scala 102:19]
    .io_x1(m_445_io_x1),
    .io_x2(m_445_io_x2),
    .io_x3(m_445_io_x3),
    .io_s(m_445_io_s),
    .io_cout(m_445_io_cout)
  );
  Adder m_446 ( // @[MUL.scala 102:19]
    .io_x1(m_446_io_x1),
    .io_x2(m_446_io_x2),
    .io_x3(m_446_io_x3),
    .io_s(m_446_io_s),
    .io_cout(m_446_io_cout)
  );
  Adder m_447 ( // @[MUL.scala 102:19]
    .io_x1(m_447_io_x1),
    .io_x2(m_447_io_x2),
    .io_x3(m_447_io_x3),
    .io_s(m_447_io_s),
    .io_cout(m_447_io_cout)
  );
  Adder m_448 ( // @[MUL.scala 102:19]
    .io_x1(m_448_io_x1),
    .io_x2(m_448_io_x2),
    .io_x3(m_448_io_x3),
    .io_s(m_448_io_s),
    .io_cout(m_448_io_cout)
  );
  Adder m_449 ( // @[MUL.scala 102:19]
    .io_x1(m_449_io_x1),
    .io_x2(m_449_io_x2),
    .io_x3(m_449_io_x3),
    .io_s(m_449_io_s),
    .io_cout(m_449_io_cout)
  );
  Adder m_450 ( // @[MUL.scala 102:19]
    .io_x1(m_450_io_x1),
    .io_x2(m_450_io_x2),
    .io_x3(m_450_io_x3),
    .io_s(m_450_io_s),
    .io_cout(m_450_io_cout)
  );
  Adder m_451 ( // @[MUL.scala 102:19]
    .io_x1(m_451_io_x1),
    .io_x2(m_451_io_x2),
    .io_x3(m_451_io_x3),
    .io_s(m_451_io_s),
    .io_cout(m_451_io_cout)
  );
  Adder m_452 ( // @[MUL.scala 102:19]
    .io_x1(m_452_io_x1),
    .io_x2(m_452_io_x2),
    .io_x3(m_452_io_x3),
    .io_s(m_452_io_s),
    .io_cout(m_452_io_cout)
  );
  Adder m_453 ( // @[MUL.scala 102:19]
    .io_x1(m_453_io_x1),
    .io_x2(m_453_io_x2),
    .io_x3(m_453_io_x3),
    .io_s(m_453_io_s),
    .io_cout(m_453_io_cout)
  );
  Adder m_454 ( // @[MUL.scala 102:19]
    .io_x1(m_454_io_x1),
    .io_x2(m_454_io_x2),
    .io_x3(m_454_io_x3),
    .io_s(m_454_io_s),
    .io_cout(m_454_io_cout)
  );
  Adder m_455 ( // @[MUL.scala 102:19]
    .io_x1(m_455_io_x1),
    .io_x2(m_455_io_x2),
    .io_x3(m_455_io_x3),
    .io_s(m_455_io_s),
    .io_cout(m_455_io_cout)
  );
  Adder m_456 ( // @[MUL.scala 102:19]
    .io_x1(m_456_io_x1),
    .io_x2(m_456_io_x2),
    .io_x3(m_456_io_x3),
    .io_s(m_456_io_s),
    .io_cout(m_456_io_cout)
  );
  Adder m_457 ( // @[MUL.scala 102:19]
    .io_x1(m_457_io_x1),
    .io_x2(m_457_io_x2),
    .io_x3(m_457_io_x3),
    .io_s(m_457_io_s),
    .io_cout(m_457_io_cout)
  );
  Adder m_458 ( // @[MUL.scala 102:19]
    .io_x1(m_458_io_x1),
    .io_x2(m_458_io_x2),
    .io_x3(m_458_io_x3),
    .io_s(m_458_io_s),
    .io_cout(m_458_io_cout)
  );
  Adder m_459 ( // @[MUL.scala 102:19]
    .io_x1(m_459_io_x1),
    .io_x2(m_459_io_x2),
    .io_x3(m_459_io_x3),
    .io_s(m_459_io_s),
    .io_cout(m_459_io_cout)
  );
  Adder m_460 ( // @[MUL.scala 102:19]
    .io_x1(m_460_io_x1),
    .io_x2(m_460_io_x2),
    .io_x3(m_460_io_x3),
    .io_s(m_460_io_s),
    .io_cout(m_460_io_cout)
  );
  Adder m_461 ( // @[MUL.scala 102:19]
    .io_x1(m_461_io_x1),
    .io_x2(m_461_io_x2),
    .io_x3(m_461_io_x3),
    .io_s(m_461_io_s),
    .io_cout(m_461_io_cout)
  );
  Adder m_462 ( // @[MUL.scala 102:19]
    .io_x1(m_462_io_x1),
    .io_x2(m_462_io_x2),
    .io_x3(m_462_io_x3),
    .io_s(m_462_io_s),
    .io_cout(m_462_io_cout)
  );
  Adder m_463 ( // @[MUL.scala 102:19]
    .io_x1(m_463_io_x1),
    .io_x2(m_463_io_x2),
    .io_x3(m_463_io_x3),
    .io_s(m_463_io_s),
    .io_cout(m_463_io_cout)
  );
  Adder m_464 ( // @[MUL.scala 102:19]
    .io_x1(m_464_io_x1),
    .io_x2(m_464_io_x2),
    .io_x3(m_464_io_x3),
    .io_s(m_464_io_s),
    .io_cout(m_464_io_cout)
  );
  Adder m_465 ( // @[MUL.scala 102:19]
    .io_x1(m_465_io_x1),
    .io_x2(m_465_io_x2),
    .io_x3(m_465_io_x3),
    .io_s(m_465_io_s),
    .io_cout(m_465_io_cout)
  );
  Adder m_466 ( // @[MUL.scala 102:19]
    .io_x1(m_466_io_x1),
    .io_x2(m_466_io_x2),
    .io_x3(m_466_io_x3),
    .io_s(m_466_io_s),
    .io_cout(m_466_io_cout)
  );
  Adder m_467 ( // @[MUL.scala 102:19]
    .io_x1(m_467_io_x1),
    .io_x2(m_467_io_x2),
    .io_x3(m_467_io_x3),
    .io_s(m_467_io_s),
    .io_cout(m_467_io_cout)
  );
  Adder m_468 ( // @[MUL.scala 102:19]
    .io_x1(m_468_io_x1),
    .io_x2(m_468_io_x2),
    .io_x3(m_468_io_x3),
    .io_s(m_468_io_s),
    .io_cout(m_468_io_cout)
  );
  Adder m_469 ( // @[MUL.scala 102:19]
    .io_x1(m_469_io_x1),
    .io_x2(m_469_io_x2),
    .io_x3(m_469_io_x3),
    .io_s(m_469_io_s),
    .io_cout(m_469_io_cout)
  );
  Adder m_470 ( // @[MUL.scala 102:19]
    .io_x1(m_470_io_x1),
    .io_x2(m_470_io_x2),
    .io_x3(m_470_io_x3),
    .io_s(m_470_io_s),
    .io_cout(m_470_io_cout)
  );
  Adder m_471 ( // @[MUL.scala 102:19]
    .io_x1(m_471_io_x1),
    .io_x2(m_471_io_x2),
    .io_x3(m_471_io_x3),
    .io_s(m_471_io_s),
    .io_cout(m_471_io_cout)
  );
  Half_Adder m_472 ( // @[MUL.scala 124:19]
    .io_in_0(m_472_io_in_0),
    .io_in_1(m_472_io_in_1),
    .io_out_0(m_472_io_out_0),
    .io_out_1(m_472_io_out_1)
  );
  Adder m_473 ( // @[MUL.scala 102:19]
    .io_x1(m_473_io_x1),
    .io_x2(m_473_io_x2),
    .io_x3(m_473_io_x3),
    .io_s(m_473_io_s),
    .io_cout(m_473_io_cout)
  );
  Adder m_474 ( // @[MUL.scala 102:19]
    .io_x1(m_474_io_x1),
    .io_x2(m_474_io_x2),
    .io_x3(m_474_io_x3),
    .io_s(m_474_io_s),
    .io_cout(m_474_io_cout)
  );
  Adder m_475 ( // @[MUL.scala 102:19]
    .io_x1(m_475_io_x1),
    .io_x2(m_475_io_x2),
    .io_x3(m_475_io_x3),
    .io_s(m_475_io_s),
    .io_cout(m_475_io_cout)
  );
  Adder m_476 ( // @[MUL.scala 102:19]
    .io_x1(m_476_io_x1),
    .io_x2(m_476_io_x2),
    .io_x3(m_476_io_x3),
    .io_s(m_476_io_s),
    .io_cout(m_476_io_cout)
  );
  Adder m_477 ( // @[MUL.scala 102:19]
    .io_x1(m_477_io_x1),
    .io_x2(m_477_io_x2),
    .io_x3(m_477_io_x3),
    .io_s(m_477_io_s),
    .io_cout(m_477_io_cout)
  );
  Adder m_478 ( // @[MUL.scala 102:19]
    .io_x1(m_478_io_x1),
    .io_x2(m_478_io_x2),
    .io_x3(m_478_io_x3),
    .io_s(m_478_io_s),
    .io_cout(m_478_io_cout)
  );
  Adder m_479 ( // @[MUL.scala 102:19]
    .io_x1(m_479_io_x1),
    .io_x2(m_479_io_x2),
    .io_x3(m_479_io_x3),
    .io_s(m_479_io_s),
    .io_cout(m_479_io_cout)
  );
  Adder m_480 ( // @[MUL.scala 102:19]
    .io_x1(m_480_io_x1),
    .io_x2(m_480_io_x2),
    .io_x3(m_480_io_x3),
    .io_s(m_480_io_s),
    .io_cout(m_480_io_cout)
  );
  Adder m_481 ( // @[MUL.scala 102:19]
    .io_x1(m_481_io_x1),
    .io_x2(m_481_io_x2),
    .io_x3(m_481_io_x3),
    .io_s(m_481_io_s),
    .io_cout(m_481_io_cout)
  );
  Adder m_482 ( // @[MUL.scala 102:19]
    .io_x1(m_482_io_x1),
    .io_x2(m_482_io_x2),
    .io_x3(m_482_io_x3),
    .io_s(m_482_io_s),
    .io_cout(m_482_io_cout)
  );
  Adder m_483 ( // @[MUL.scala 102:19]
    .io_x1(m_483_io_x1),
    .io_x2(m_483_io_x2),
    .io_x3(m_483_io_x3),
    .io_s(m_483_io_s),
    .io_cout(m_483_io_cout)
  );
  Adder m_484 ( // @[MUL.scala 102:19]
    .io_x1(m_484_io_x1),
    .io_x2(m_484_io_x2),
    .io_x3(m_484_io_x3),
    .io_s(m_484_io_s),
    .io_cout(m_484_io_cout)
  );
  Adder m_485 ( // @[MUL.scala 102:19]
    .io_x1(m_485_io_x1),
    .io_x2(m_485_io_x2),
    .io_x3(m_485_io_x3),
    .io_s(m_485_io_s),
    .io_cout(m_485_io_cout)
  );
  Adder m_486 ( // @[MUL.scala 102:19]
    .io_x1(m_486_io_x1),
    .io_x2(m_486_io_x2),
    .io_x3(m_486_io_x3),
    .io_s(m_486_io_s),
    .io_cout(m_486_io_cout)
  );
  Adder m_487 ( // @[MUL.scala 102:19]
    .io_x1(m_487_io_x1),
    .io_x2(m_487_io_x2),
    .io_x3(m_487_io_x3),
    .io_s(m_487_io_s),
    .io_cout(m_487_io_cout)
  );
  Adder m_488 ( // @[MUL.scala 102:19]
    .io_x1(m_488_io_x1),
    .io_x2(m_488_io_x2),
    .io_x3(m_488_io_x3),
    .io_s(m_488_io_s),
    .io_cout(m_488_io_cout)
  );
  Adder m_489 ( // @[MUL.scala 102:19]
    .io_x1(m_489_io_x1),
    .io_x2(m_489_io_x2),
    .io_x3(m_489_io_x3),
    .io_s(m_489_io_s),
    .io_cout(m_489_io_cout)
  );
  Adder m_490 ( // @[MUL.scala 102:19]
    .io_x1(m_490_io_x1),
    .io_x2(m_490_io_x2),
    .io_x3(m_490_io_x3),
    .io_s(m_490_io_s),
    .io_cout(m_490_io_cout)
  );
  Adder m_491 ( // @[MUL.scala 102:19]
    .io_x1(m_491_io_x1),
    .io_x2(m_491_io_x2),
    .io_x3(m_491_io_x3),
    .io_s(m_491_io_s),
    .io_cout(m_491_io_cout)
  );
  Adder m_492 ( // @[MUL.scala 102:19]
    .io_x1(m_492_io_x1),
    .io_x2(m_492_io_x2),
    .io_x3(m_492_io_x3),
    .io_s(m_492_io_s),
    .io_cout(m_492_io_cout)
  );
  Adder m_493 ( // @[MUL.scala 102:19]
    .io_x1(m_493_io_x1),
    .io_x2(m_493_io_x2),
    .io_x3(m_493_io_x3),
    .io_s(m_493_io_s),
    .io_cout(m_493_io_cout)
  );
  Adder m_494 ( // @[MUL.scala 102:19]
    .io_x1(m_494_io_x1),
    .io_x2(m_494_io_x2),
    .io_x3(m_494_io_x3),
    .io_s(m_494_io_s),
    .io_cout(m_494_io_cout)
  );
  Adder m_495 ( // @[MUL.scala 102:19]
    .io_x1(m_495_io_x1),
    .io_x2(m_495_io_x2),
    .io_x3(m_495_io_x3),
    .io_s(m_495_io_s),
    .io_cout(m_495_io_cout)
  );
  Adder m_496 ( // @[MUL.scala 102:19]
    .io_x1(m_496_io_x1),
    .io_x2(m_496_io_x2),
    .io_x3(m_496_io_x3),
    .io_s(m_496_io_s),
    .io_cout(m_496_io_cout)
  );
  Adder m_497 ( // @[MUL.scala 102:19]
    .io_x1(m_497_io_x1),
    .io_x2(m_497_io_x2),
    .io_x3(m_497_io_x3),
    .io_s(m_497_io_s),
    .io_cout(m_497_io_cout)
  );
  Adder m_498 ( // @[MUL.scala 102:19]
    .io_x1(m_498_io_x1),
    .io_x2(m_498_io_x2),
    .io_x3(m_498_io_x3),
    .io_s(m_498_io_s),
    .io_cout(m_498_io_cout)
  );
  Adder m_499 ( // @[MUL.scala 102:19]
    .io_x1(m_499_io_x1),
    .io_x2(m_499_io_x2),
    .io_x3(m_499_io_x3),
    .io_s(m_499_io_s),
    .io_cout(m_499_io_cout)
  );
  Adder m_500 ( // @[MUL.scala 102:19]
    .io_x1(m_500_io_x1),
    .io_x2(m_500_io_x2),
    .io_x3(m_500_io_x3),
    .io_s(m_500_io_s),
    .io_cout(m_500_io_cout)
  );
  Adder m_501 ( // @[MUL.scala 102:19]
    .io_x1(m_501_io_x1),
    .io_x2(m_501_io_x2),
    .io_x3(m_501_io_x3),
    .io_s(m_501_io_s),
    .io_cout(m_501_io_cout)
  );
  Adder m_502 ( // @[MUL.scala 102:19]
    .io_x1(m_502_io_x1),
    .io_x2(m_502_io_x2),
    .io_x3(m_502_io_x3),
    .io_s(m_502_io_s),
    .io_cout(m_502_io_cout)
  );
  Adder m_503 ( // @[MUL.scala 102:19]
    .io_x1(m_503_io_x1),
    .io_x2(m_503_io_x2),
    .io_x3(m_503_io_x3),
    .io_s(m_503_io_s),
    .io_cout(m_503_io_cout)
  );
  Adder m_504 ( // @[MUL.scala 102:19]
    .io_x1(m_504_io_x1),
    .io_x2(m_504_io_x2),
    .io_x3(m_504_io_x3),
    .io_s(m_504_io_s),
    .io_cout(m_504_io_cout)
  );
  Adder m_505 ( // @[MUL.scala 102:19]
    .io_x1(m_505_io_x1),
    .io_x2(m_505_io_x2),
    .io_x3(m_505_io_x3),
    .io_s(m_505_io_s),
    .io_cout(m_505_io_cout)
  );
  Adder m_506 ( // @[MUL.scala 102:19]
    .io_x1(m_506_io_x1),
    .io_x2(m_506_io_x2),
    .io_x3(m_506_io_x3),
    .io_s(m_506_io_s),
    .io_cout(m_506_io_cout)
  );
  Adder m_507 ( // @[MUL.scala 102:19]
    .io_x1(m_507_io_x1),
    .io_x2(m_507_io_x2),
    .io_x3(m_507_io_x3),
    .io_s(m_507_io_s),
    .io_cout(m_507_io_cout)
  );
  Adder m_508 ( // @[MUL.scala 102:19]
    .io_x1(m_508_io_x1),
    .io_x2(m_508_io_x2),
    .io_x3(m_508_io_x3),
    .io_s(m_508_io_s),
    .io_cout(m_508_io_cout)
  );
  Adder m_509 ( // @[MUL.scala 102:19]
    .io_x1(m_509_io_x1),
    .io_x2(m_509_io_x2),
    .io_x3(m_509_io_x3),
    .io_s(m_509_io_s),
    .io_cout(m_509_io_cout)
  );
  Adder m_510 ( // @[MUL.scala 102:19]
    .io_x1(m_510_io_x1),
    .io_x2(m_510_io_x2),
    .io_x3(m_510_io_x3),
    .io_s(m_510_io_s),
    .io_cout(m_510_io_cout)
  );
  Adder m_511 ( // @[MUL.scala 102:19]
    .io_x1(m_511_io_x1),
    .io_x2(m_511_io_x2),
    .io_x3(m_511_io_x3),
    .io_s(m_511_io_s),
    .io_cout(m_511_io_cout)
  );
  Adder m_512 ( // @[MUL.scala 102:19]
    .io_x1(m_512_io_x1),
    .io_x2(m_512_io_x2),
    .io_x3(m_512_io_x3),
    .io_s(m_512_io_s),
    .io_cout(m_512_io_cout)
  );
  Adder m_513 ( // @[MUL.scala 102:19]
    .io_x1(m_513_io_x1),
    .io_x2(m_513_io_x2),
    .io_x3(m_513_io_x3),
    .io_s(m_513_io_s),
    .io_cout(m_513_io_cout)
  );
  Adder m_514 ( // @[MUL.scala 102:19]
    .io_x1(m_514_io_x1),
    .io_x2(m_514_io_x2),
    .io_x3(m_514_io_x3),
    .io_s(m_514_io_s),
    .io_cout(m_514_io_cout)
  );
  Adder m_515 ( // @[MUL.scala 102:19]
    .io_x1(m_515_io_x1),
    .io_x2(m_515_io_x2),
    .io_x3(m_515_io_x3),
    .io_s(m_515_io_s),
    .io_cout(m_515_io_cout)
  );
  Adder m_516 ( // @[MUL.scala 102:19]
    .io_x1(m_516_io_x1),
    .io_x2(m_516_io_x2),
    .io_x3(m_516_io_x3),
    .io_s(m_516_io_s),
    .io_cout(m_516_io_cout)
  );
  Adder m_517 ( // @[MUL.scala 102:19]
    .io_x1(m_517_io_x1),
    .io_x2(m_517_io_x2),
    .io_x3(m_517_io_x3),
    .io_s(m_517_io_s),
    .io_cout(m_517_io_cout)
  );
  Adder m_518 ( // @[MUL.scala 102:19]
    .io_x1(m_518_io_x1),
    .io_x2(m_518_io_x2),
    .io_x3(m_518_io_x3),
    .io_s(m_518_io_s),
    .io_cout(m_518_io_cout)
  );
  Adder m_519 ( // @[MUL.scala 102:19]
    .io_x1(m_519_io_x1),
    .io_x2(m_519_io_x2),
    .io_x3(m_519_io_x3),
    .io_s(m_519_io_s),
    .io_cout(m_519_io_cout)
  );
  Adder m_520 ( // @[MUL.scala 102:19]
    .io_x1(m_520_io_x1),
    .io_x2(m_520_io_x2),
    .io_x3(m_520_io_x3),
    .io_s(m_520_io_s),
    .io_cout(m_520_io_cout)
  );
  Adder m_521 ( // @[MUL.scala 102:19]
    .io_x1(m_521_io_x1),
    .io_x2(m_521_io_x2),
    .io_x3(m_521_io_x3),
    .io_s(m_521_io_s),
    .io_cout(m_521_io_cout)
  );
  Half_Adder m_522 ( // @[MUL.scala 124:19]
    .io_in_0(m_522_io_in_0),
    .io_in_1(m_522_io_in_1),
    .io_out_0(m_522_io_out_0),
    .io_out_1(m_522_io_out_1)
  );
  Adder m_523 ( // @[MUL.scala 102:19]
    .io_x1(m_523_io_x1),
    .io_x2(m_523_io_x2),
    .io_x3(m_523_io_x3),
    .io_s(m_523_io_s),
    .io_cout(m_523_io_cout)
  );
  Adder m_524 ( // @[MUL.scala 102:19]
    .io_x1(m_524_io_x1),
    .io_x2(m_524_io_x2),
    .io_x3(m_524_io_x3),
    .io_s(m_524_io_s),
    .io_cout(m_524_io_cout)
  );
  Adder m_525 ( // @[MUL.scala 102:19]
    .io_x1(m_525_io_x1),
    .io_x2(m_525_io_x2),
    .io_x3(m_525_io_x3),
    .io_s(m_525_io_s),
    .io_cout(m_525_io_cout)
  );
  Adder m_526 ( // @[MUL.scala 102:19]
    .io_x1(m_526_io_x1),
    .io_x2(m_526_io_x2),
    .io_x3(m_526_io_x3),
    .io_s(m_526_io_s),
    .io_cout(m_526_io_cout)
  );
  Adder m_527 ( // @[MUL.scala 102:19]
    .io_x1(m_527_io_x1),
    .io_x2(m_527_io_x2),
    .io_x3(m_527_io_x3),
    .io_s(m_527_io_s),
    .io_cout(m_527_io_cout)
  );
  Adder m_528 ( // @[MUL.scala 102:19]
    .io_x1(m_528_io_x1),
    .io_x2(m_528_io_x2),
    .io_x3(m_528_io_x3),
    .io_s(m_528_io_s),
    .io_cout(m_528_io_cout)
  );
  Adder m_529 ( // @[MUL.scala 102:19]
    .io_x1(m_529_io_x1),
    .io_x2(m_529_io_x2),
    .io_x3(m_529_io_x3),
    .io_s(m_529_io_s),
    .io_cout(m_529_io_cout)
  );
  Adder m_530 ( // @[MUL.scala 102:19]
    .io_x1(m_530_io_x1),
    .io_x2(m_530_io_x2),
    .io_x3(m_530_io_x3),
    .io_s(m_530_io_s),
    .io_cout(m_530_io_cout)
  );
  Adder m_531 ( // @[MUL.scala 102:19]
    .io_x1(m_531_io_x1),
    .io_x2(m_531_io_x2),
    .io_x3(m_531_io_x3),
    .io_s(m_531_io_s),
    .io_cout(m_531_io_cout)
  );
  Half_Adder m_532 ( // @[MUL.scala 124:19]
    .io_in_0(m_532_io_in_0),
    .io_in_1(m_532_io_in_1),
    .io_out_0(m_532_io_out_0),
    .io_out_1(m_532_io_out_1)
  );
  Adder m_533 ( // @[MUL.scala 102:19]
    .io_x1(m_533_io_x1),
    .io_x2(m_533_io_x2),
    .io_x3(m_533_io_x3),
    .io_s(m_533_io_s),
    .io_cout(m_533_io_cout)
  );
  Adder m_534 ( // @[MUL.scala 102:19]
    .io_x1(m_534_io_x1),
    .io_x2(m_534_io_x2),
    .io_x3(m_534_io_x3),
    .io_s(m_534_io_s),
    .io_cout(m_534_io_cout)
  );
  Adder m_535 ( // @[MUL.scala 102:19]
    .io_x1(m_535_io_x1),
    .io_x2(m_535_io_x2),
    .io_x3(m_535_io_x3),
    .io_s(m_535_io_s),
    .io_cout(m_535_io_cout)
  );
  Adder m_536 ( // @[MUL.scala 102:19]
    .io_x1(m_536_io_x1),
    .io_x2(m_536_io_x2),
    .io_x3(m_536_io_x3),
    .io_s(m_536_io_s),
    .io_cout(m_536_io_cout)
  );
  Adder m_537 ( // @[MUL.scala 102:19]
    .io_x1(m_537_io_x1),
    .io_x2(m_537_io_x2),
    .io_x3(m_537_io_x3),
    .io_s(m_537_io_s),
    .io_cout(m_537_io_cout)
  );
  Adder m_538 ( // @[MUL.scala 102:19]
    .io_x1(m_538_io_x1),
    .io_x2(m_538_io_x2),
    .io_x3(m_538_io_x3),
    .io_s(m_538_io_s),
    .io_cout(m_538_io_cout)
  );
  Adder m_539 ( // @[MUL.scala 102:19]
    .io_x1(m_539_io_x1),
    .io_x2(m_539_io_x2),
    .io_x3(m_539_io_x3),
    .io_s(m_539_io_s),
    .io_cout(m_539_io_cout)
  );
  Adder m_540 ( // @[MUL.scala 102:19]
    .io_x1(m_540_io_x1),
    .io_x2(m_540_io_x2),
    .io_x3(m_540_io_x3),
    .io_s(m_540_io_s),
    .io_cout(m_540_io_cout)
  );
  Adder m_541 ( // @[MUL.scala 102:19]
    .io_x1(m_541_io_x1),
    .io_x2(m_541_io_x2),
    .io_x3(m_541_io_x3),
    .io_s(m_541_io_s),
    .io_cout(m_541_io_cout)
  );
  Adder m_542 ( // @[MUL.scala 102:19]
    .io_x1(m_542_io_x1),
    .io_x2(m_542_io_x2),
    .io_x3(m_542_io_x3),
    .io_s(m_542_io_s),
    .io_cout(m_542_io_cout)
  );
  Adder m_543 ( // @[MUL.scala 102:19]
    .io_x1(m_543_io_x1),
    .io_x2(m_543_io_x2),
    .io_x3(m_543_io_x3),
    .io_s(m_543_io_s),
    .io_cout(m_543_io_cout)
  );
  Adder m_544 ( // @[MUL.scala 102:19]
    .io_x1(m_544_io_x1),
    .io_x2(m_544_io_x2),
    .io_x3(m_544_io_x3),
    .io_s(m_544_io_s),
    .io_cout(m_544_io_cout)
  );
  Adder m_545 ( // @[MUL.scala 102:19]
    .io_x1(m_545_io_x1),
    .io_x2(m_545_io_x2),
    .io_x3(m_545_io_x3),
    .io_s(m_545_io_s),
    .io_cout(m_545_io_cout)
  );
  Adder m_546 ( // @[MUL.scala 102:19]
    .io_x1(m_546_io_x1),
    .io_x2(m_546_io_x2),
    .io_x3(m_546_io_x3),
    .io_s(m_546_io_s),
    .io_cout(m_546_io_cout)
  );
  Adder m_547 ( // @[MUL.scala 102:19]
    .io_x1(m_547_io_x1),
    .io_x2(m_547_io_x2),
    .io_x3(m_547_io_x3),
    .io_s(m_547_io_s),
    .io_cout(m_547_io_cout)
  );
  Adder m_548 ( // @[MUL.scala 102:19]
    .io_x1(m_548_io_x1),
    .io_x2(m_548_io_x2),
    .io_x3(m_548_io_x3),
    .io_s(m_548_io_s),
    .io_cout(m_548_io_cout)
  );
  Adder m_549 ( // @[MUL.scala 102:19]
    .io_x1(m_549_io_x1),
    .io_x2(m_549_io_x2),
    .io_x3(m_549_io_x3),
    .io_s(m_549_io_s),
    .io_cout(m_549_io_cout)
  );
  Adder m_550 ( // @[MUL.scala 102:19]
    .io_x1(m_550_io_x1),
    .io_x2(m_550_io_x2),
    .io_x3(m_550_io_x3),
    .io_s(m_550_io_s),
    .io_cout(m_550_io_cout)
  );
  Adder m_551 ( // @[MUL.scala 102:19]
    .io_x1(m_551_io_x1),
    .io_x2(m_551_io_x2),
    .io_x3(m_551_io_x3),
    .io_s(m_551_io_s),
    .io_cout(m_551_io_cout)
  );
  Adder m_552 ( // @[MUL.scala 102:19]
    .io_x1(m_552_io_x1),
    .io_x2(m_552_io_x2),
    .io_x3(m_552_io_x3),
    .io_s(m_552_io_s),
    .io_cout(m_552_io_cout)
  );
  Adder m_553 ( // @[MUL.scala 102:19]
    .io_x1(m_553_io_x1),
    .io_x2(m_553_io_x2),
    .io_x3(m_553_io_x3),
    .io_s(m_553_io_s),
    .io_cout(m_553_io_cout)
  );
  Adder m_554 ( // @[MUL.scala 102:19]
    .io_x1(m_554_io_x1),
    .io_x2(m_554_io_x2),
    .io_x3(m_554_io_x3),
    .io_s(m_554_io_s),
    .io_cout(m_554_io_cout)
  );
  Adder m_555 ( // @[MUL.scala 102:19]
    .io_x1(m_555_io_x1),
    .io_x2(m_555_io_x2),
    .io_x3(m_555_io_x3),
    .io_s(m_555_io_s),
    .io_cout(m_555_io_cout)
  );
  Adder m_556 ( // @[MUL.scala 102:19]
    .io_x1(m_556_io_x1),
    .io_x2(m_556_io_x2),
    .io_x3(m_556_io_x3),
    .io_s(m_556_io_s),
    .io_cout(m_556_io_cout)
  );
  Adder m_557 ( // @[MUL.scala 102:19]
    .io_x1(m_557_io_x1),
    .io_x2(m_557_io_x2),
    .io_x3(m_557_io_x3),
    .io_s(m_557_io_s),
    .io_cout(m_557_io_cout)
  );
  Adder m_558 ( // @[MUL.scala 102:19]
    .io_x1(m_558_io_x1),
    .io_x2(m_558_io_x2),
    .io_x3(m_558_io_x3),
    .io_s(m_558_io_s),
    .io_cout(m_558_io_cout)
  );
  Adder m_559 ( // @[MUL.scala 102:19]
    .io_x1(m_559_io_x1),
    .io_x2(m_559_io_x2),
    .io_x3(m_559_io_x3),
    .io_s(m_559_io_s),
    .io_cout(m_559_io_cout)
  );
  Adder m_560 ( // @[MUL.scala 102:19]
    .io_x1(m_560_io_x1),
    .io_x2(m_560_io_x2),
    .io_x3(m_560_io_x3),
    .io_s(m_560_io_s),
    .io_cout(m_560_io_cout)
  );
  Adder m_561 ( // @[MUL.scala 102:19]
    .io_x1(m_561_io_x1),
    .io_x2(m_561_io_x2),
    .io_x3(m_561_io_x3),
    .io_s(m_561_io_s),
    .io_cout(m_561_io_cout)
  );
  Adder m_562 ( // @[MUL.scala 102:19]
    .io_x1(m_562_io_x1),
    .io_x2(m_562_io_x2),
    .io_x3(m_562_io_x3),
    .io_s(m_562_io_s),
    .io_cout(m_562_io_cout)
  );
  Adder m_563 ( // @[MUL.scala 102:19]
    .io_x1(m_563_io_x1),
    .io_x2(m_563_io_x2),
    .io_x3(m_563_io_x3),
    .io_s(m_563_io_s),
    .io_cout(m_563_io_cout)
  );
  Adder m_564 ( // @[MUL.scala 102:19]
    .io_x1(m_564_io_x1),
    .io_x2(m_564_io_x2),
    .io_x3(m_564_io_x3),
    .io_s(m_564_io_s),
    .io_cout(m_564_io_cout)
  );
  Adder m_565 ( // @[MUL.scala 102:19]
    .io_x1(m_565_io_x1),
    .io_x2(m_565_io_x2),
    .io_x3(m_565_io_x3),
    .io_s(m_565_io_s),
    .io_cout(m_565_io_cout)
  );
  Adder m_566 ( // @[MUL.scala 102:19]
    .io_x1(m_566_io_x1),
    .io_x2(m_566_io_x2),
    .io_x3(m_566_io_x3),
    .io_s(m_566_io_s),
    .io_cout(m_566_io_cout)
  );
  Adder m_567 ( // @[MUL.scala 102:19]
    .io_x1(m_567_io_x1),
    .io_x2(m_567_io_x2),
    .io_x3(m_567_io_x3),
    .io_s(m_567_io_s),
    .io_cout(m_567_io_cout)
  );
  Adder m_568 ( // @[MUL.scala 102:19]
    .io_x1(m_568_io_x1),
    .io_x2(m_568_io_x2),
    .io_x3(m_568_io_x3),
    .io_s(m_568_io_s),
    .io_cout(m_568_io_cout)
  );
  Adder m_569 ( // @[MUL.scala 102:19]
    .io_x1(m_569_io_x1),
    .io_x2(m_569_io_x2),
    .io_x3(m_569_io_x3),
    .io_s(m_569_io_s),
    .io_cout(m_569_io_cout)
  );
  Adder m_570 ( // @[MUL.scala 102:19]
    .io_x1(m_570_io_x1),
    .io_x2(m_570_io_x2),
    .io_x3(m_570_io_x3),
    .io_s(m_570_io_s),
    .io_cout(m_570_io_cout)
  );
  Adder m_571 ( // @[MUL.scala 102:19]
    .io_x1(m_571_io_x1),
    .io_x2(m_571_io_x2),
    .io_x3(m_571_io_x3),
    .io_s(m_571_io_s),
    .io_cout(m_571_io_cout)
  );
  Adder m_572 ( // @[MUL.scala 102:19]
    .io_x1(m_572_io_x1),
    .io_x2(m_572_io_x2),
    .io_x3(m_572_io_x3),
    .io_s(m_572_io_s),
    .io_cout(m_572_io_cout)
  );
  Adder m_573 ( // @[MUL.scala 102:19]
    .io_x1(m_573_io_x1),
    .io_x2(m_573_io_x2),
    .io_x3(m_573_io_x3),
    .io_s(m_573_io_s),
    .io_cout(m_573_io_cout)
  );
  Adder m_574 ( // @[MUL.scala 102:19]
    .io_x1(m_574_io_x1),
    .io_x2(m_574_io_x2),
    .io_x3(m_574_io_x3),
    .io_s(m_574_io_s),
    .io_cout(m_574_io_cout)
  );
  Adder m_575 ( // @[MUL.scala 102:19]
    .io_x1(m_575_io_x1),
    .io_x2(m_575_io_x2),
    .io_x3(m_575_io_x3),
    .io_s(m_575_io_s),
    .io_cout(m_575_io_cout)
  );
  Adder m_576 ( // @[MUL.scala 102:19]
    .io_x1(m_576_io_x1),
    .io_x2(m_576_io_x2),
    .io_x3(m_576_io_x3),
    .io_s(m_576_io_s),
    .io_cout(m_576_io_cout)
  );
  Half_Adder m_577 ( // @[MUL.scala 124:19]
    .io_in_0(m_577_io_in_0),
    .io_in_1(m_577_io_in_1),
    .io_out_0(m_577_io_out_0),
    .io_out_1(m_577_io_out_1)
  );
  Adder m_578 ( // @[MUL.scala 102:19]
    .io_x1(m_578_io_x1),
    .io_x2(m_578_io_x2),
    .io_x3(m_578_io_x3),
    .io_s(m_578_io_s),
    .io_cout(m_578_io_cout)
  );
  Adder m_579 ( // @[MUL.scala 102:19]
    .io_x1(m_579_io_x1),
    .io_x2(m_579_io_x2),
    .io_x3(m_579_io_x3),
    .io_s(m_579_io_s),
    .io_cout(m_579_io_cout)
  );
  Adder m_580 ( // @[MUL.scala 102:19]
    .io_x1(m_580_io_x1),
    .io_x2(m_580_io_x2),
    .io_x3(m_580_io_x3),
    .io_s(m_580_io_s),
    .io_cout(m_580_io_cout)
  );
  Adder m_581 ( // @[MUL.scala 102:19]
    .io_x1(m_581_io_x1),
    .io_x2(m_581_io_x2),
    .io_x3(m_581_io_x3),
    .io_s(m_581_io_s),
    .io_cout(m_581_io_cout)
  );
  Adder m_582 ( // @[MUL.scala 102:19]
    .io_x1(m_582_io_x1),
    .io_x2(m_582_io_x2),
    .io_x3(m_582_io_x3),
    .io_s(m_582_io_s),
    .io_cout(m_582_io_cout)
  );
  Adder m_583 ( // @[MUL.scala 102:19]
    .io_x1(m_583_io_x1),
    .io_x2(m_583_io_x2),
    .io_x3(m_583_io_x3),
    .io_s(m_583_io_s),
    .io_cout(m_583_io_cout)
  );
  Adder m_584 ( // @[MUL.scala 102:19]
    .io_x1(m_584_io_x1),
    .io_x2(m_584_io_x2),
    .io_x3(m_584_io_x3),
    .io_s(m_584_io_s),
    .io_cout(m_584_io_cout)
  );
  Adder m_585 ( // @[MUL.scala 102:19]
    .io_x1(m_585_io_x1),
    .io_x2(m_585_io_x2),
    .io_x3(m_585_io_x3),
    .io_s(m_585_io_s),
    .io_cout(m_585_io_cout)
  );
  Half_Adder m_586 ( // @[MUL.scala 124:19]
    .io_in_0(m_586_io_in_0),
    .io_in_1(m_586_io_in_1),
    .io_out_0(m_586_io_out_0),
    .io_out_1(m_586_io_out_1)
  );
  Adder m_587 ( // @[MUL.scala 102:19]
    .io_x1(m_587_io_x1),
    .io_x2(m_587_io_x2),
    .io_x3(m_587_io_x3),
    .io_s(m_587_io_s),
    .io_cout(m_587_io_cout)
  );
  Adder m_588 ( // @[MUL.scala 102:19]
    .io_x1(m_588_io_x1),
    .io_x2(m_588_io_x2),
    .io_x3(m_588_io_x3),
    .io_s(m_588_io_s),
    .io_cout(m_588_io_cout)
  );
  Adder m_589 ( // @[MUL.scala 102:19]
    .io_x1(m_589_io_x1),
    .io_x2(m_589_io_x2),
    .io_x3(m_589_io_x3),
    .io_s(m_589_io_s),
    .io_cout(m_589_io_cout)
  );
  Adder m_590 ( // @[MUL.scala 102:19]
    .io_x1(m_590_io_x1),
    .io_x2(m_590_io_x2),
    .io_x3(m_590_io_x3),
    .io_s(m_590_io_s),
    .io_cout(m_590_io_cout)
  );
  Adder m_591 ( // @[MUL.scala 102:19]
    .io_x1(m_591_io_x1),
    .io_x2(m_591_io_x2),
    .io_x3(m_591_io_x3),
    .io_s(m_591_io_s),
    .io_cout(m_591_io_cout)
  );
  Adder m_592 ( // @[MUL.scala 102:19]
    .io_x1(m_592_io_x1),
    .io_x2(m_592_io_x2),
    .io_x3(m_592_io_x3),
    .io_s(m_592_io_s),
    .io_cout(m_592_io_cout)
  );
  Adder m_593 ( // @[MUL.scala 102:19]
    .io_x1(m_593_io_x1),
    .io_x2(m_593_io_x2),
    .io_x3(m_593_io_x3),
    .io_s(m_593_io_s),
    .io_cout(m_593_io_cout)
  );
  Adder m_594 ( // @[MUL.scala 102:19]
    .io_x1(m_594_io_x1),
    .io_x2(m_594_io_x2),
    .io_x3(m_594_io_x3),
    .io_s(m_594_io_s),
    .io_cout(m_594_io_cout)
  );
  Adder m_595 ( // @[MUL.scala 102:19]
    .io_x1(m_595_io_x1),
    .io_x2(m_595_io_x2),
    .io_x3(m_595_io_x3),
    .io_s(m_595_io_s),
    .io_cout(m_595_io_cout)
  );
  Adder m_596 ( // @[MUL.scala 102:19]
    .io_x1(m_596_io_x1),
    .io_x2(m_596_io_x2),
    .io_x3(m_596_io_x3),
    .io_s(m_596_io_s),
    .io_cout(m_596_io_cout)
  );
  Adder m_597 ( // @[MUL.scala 102:19]
    .io_x1(m_597_io_x1),
    .io_x2(m_597_io_x2),
    .io_x3(m_597_io_x3),
    .io_s(m_597_io_s),
    .io_cout(m_597_io_cout)
  );
  Adder m_598 ( // @[MUL.scala 102:19]
    .io_x1(m_598_io_x1),
    .io_x2(m_598_io_x2),
    .io_x3(m_598_io_x3),
    .io_s(m_598_io_s),
    .io_cout(m_598_io_cout)
  );
  Adder m_599 ( // @[MUL.scala 102:19]
    .io_x1(m_599_io_x1),
    .io_x2(m_599_io_x2),
    .io_x3(m_599_io_x3),
    .io_s(m_599_io_s),
    .io_cout(m_599_io_cout)
  );
  Adder m_600 ( // @[MUL.scala 102:19]
    .io_x1(m_600_io_x1),
    .io_x2(m_600_io_x2),
    .io_x3(m_600_io_x3),
    .io_s(m_600_io_s),
    .io_cout(m_600_io_cout)
  );
  Adder m_601 ( // @[MUL.scala 102:19]
    .io_x1(m_601_io_x1),
    .io_x2(m_601_io_x2),
    .io_x3(m_601_io_x3),
    .io_s(m_601_io_s),
    .io_cout(m_601_io_cout)
  );
  Adder m_602 ( // @[MUL.scala 102:19]
    .io_x1(m_602_io_x1),
    .io_x2(m_602_io_x2),
    .io_x3(m_602_io_x3),
    .io_s(m_602_io_s),
    .io_cout(m_602_io_cout)
  );
  Adder m_603 ( // @[MUL.scala 102:19]
    .io_x1(m_603_io_x1),
    .io_x2(m_603_io_x2),
    .io_x3(m_603_io_x3),
    .io_s(m_603_io_s),
    .io_cout(m_603_io_cout)
  );
  Adder m_604 ( // @[MUL.scala 102:19]
    .io_x1(m_604_io_x1),
    .io_x2(m_604_io_x2),
    .io_x3(m_604_io_x3),
    .io_s(m_604_io_s),
    .io_cout(m_604_io_cout)
  );
  Adder m_605 ( // @[MUL.scala 102:19]
    .io_x1(m_605_io_x1),
    .io_x2(m_605_io_x2),
    .io_x3(m_605_io_x3),
    .io_s(m_605_io_s),
    .io_cout(m_605_io_cout)
  );
  Adder m_606 ( // @[MUL.scala 102:19]
    .io_x1(m_606_io_x1),
    .io_x2(m_606_io_x2),
    .io_x3(m_606_io_x3),
    .io_s(m_606_io_s),
    .io_cout(m_606_io_cout)
  );
  Adder m_607 ( // @[MUL.scala 102:19]
    .io_x1(m_607_io_x1),
    .io_x2(m_607_io_x2),
    .io_x3(m_607_io_x3),
    .io_s(m_607_io_s),
    .io_cout(m_607_io_cout)
  );
  Adder m_608 ( // @[MUL.scala 102:19]
    .io_x1(m_608_io_x1),
    .io_x2(m_608_io_x2),
    .io_x3(m_608_io_x3),
    .io_s(m_608_io_s),
    .io_cout(m_608_io_cout)
  );
  Adder m_609 ( // @[MUL.scala 102:19]
    .io_x1(m_609_io_x1),
    .io_x2(m_609_io_x2),
    .io_x3(m_609_io_x3),
    .io_s(m_609_io_s),
    .io_cout(m_609_io_cout)
  );
  Adder m_610 ( // @[MUL.scala 102:19]
    .io_x1(m_610_io_x1),
    .io_x2(m_610_io_x2),
    .io_x3(m_610_io_x3),
    .io_s(m_610_io_s),
    .io_cout(m_610_io_cout)
  );
  Adder m_611 ( // @[MUL.scala 102:19]
    .io_x1(m_611_io_x1),
    .io_x2(m_611_io_x2),
    .io_x3(m_611_io_x3),
    .io_s(m_611_io_s),
    .io_cout(m_611_io_cout)
  );
  Adder m_612 ( // @[MUL.scala 102:19]
    .io_x1(m_612_io_x1),
    .io_x2(m_612_io_x2),
    .io_x3(m_612_io_x3),
    .io_s(m_612_io_s),
    .io_cout(m_612_io_cout)
  );
  Adder m_613 ( // @[MUL.scala 102:19]
    .io_x1(m_613_io_x1),
    .io_x2(m_613_io_x2),
    .io_x3(m_613_io_x3),
    .io_s(m_613_io_s),
    .io_cout(m_613_io_cout)
  );
  Adder m_614 ( // @[MUL.scala 102:19]
    .io_x1(m_614_io_x1),
    .io_x2(m_614_io_x2),
    .io_x3(m_614_io_x3),
    .io_s(m_614_io_s),
    .io_cout(m_614_io_cout)
  );
  Adder m_615 ( // @[MUL.scala 102:19]
    .io_x1(m_615_io_x1),
    .io_x2(m_615_io_x2),
    .io_x3(m_615_io_x3),
    .io_s(m_615_io_s),
    .io_cout(m_615_io_cout)
  );
  Adder m_616 ( // @[MUL.scala 102:19]
    .io_x1(m_616_io_x1),
    .io_x2(m_616_io_x2),
    .io_x3(m_616_io_x3),
    .io_s(m_616_io_s),
    .io_cout(m_616_io_cout)
  );
  Adder m_617 ( // @[MUL.scala 102:19]
    .io_x1(m_617_io_x1),
    .io_x2(m_617_io_x2),
    .io_x3(m_617_io_x3),
    .io_s(m_617_io_s),
    .io_cout(m_617_io_cout)
  );
  Adder m_618 ( // @[MUL.scala 102:19]
    .io_x1(m_618_io_x1),
    .io_x2(m_618_io_x2),
    .io_x3(m_618_io_x3),
    .io_s(m_618_io_s),
    .io_cout(m_618_io_cout)
  );
  Adder m_619 ( // @[MUL.scala 102:19]
    .io_x1(m_619_io_x1),
    .io_x2(m_619_io_x2),
    .io_x3(m_619_io_x3),
    .io_s(m_619_io_s),
    .io_cout(m_619_io_cout)
  );
  Adder m_620 ( // @[MUL.scala 102:19]
    .io_x1(m_620_io_x1),
    .io_x2(m_620_io_x2),
    .io_x3(m_620_io_x3),
    .io_s(m_620_io_s),
    .io_cout(m_620_io_cout)
  );
  Adder m_621 ( // @[MUL.scala 102:19]
    .io_x1(m_621_io_x1),
    .io_x2(m_621_io_x2),
    .io_x3(m_621_io_x3),
    .io_s(m_621_io_s),
    .io_cout(m_621_io_cout)
  );
  Adder m_622 ( // @[MUL.scala 102:19]
    .io_x1(m_622_io_x1),
    .io_x2(m_622_io_x2),
    .io_x3(m_622_io_x3),
    .io_s(m_622_io_s),
    .io_cout(m_622_io_cout)
  );
  Adder m_623 ( // @[MUL.scala 102:19]
    .io_x1(m_623_io_x1),
    .io_x2(m_623_io_x2),
    .io_x3(m_623_io_x3),
    .io_s(m_623_io_s),
    .io_cout(m_623_io_cout)
  );
  Adder m_624 ( // @[MUL.scala 102:19]
    .io_x1(m_624_io_x1),
    .io_x2(m_624_io_x2),
    .io_x3(m_624_io_x3),
    .io_s(m_624_io_s),
    .io_cout(m_624_io_cout)
  );
  Adder m_625 ( // @[MUL.scala 102:19]
    .io_x1(m_625_io_x1),
    .io_x2(m_625_io_x2),
    .io_x3(m_625_io_x3),
    .io_s(m_625_io_s),
    .io_cout(m_625_io_cout)
  );
  Half_Adder m_626 ( // @[MUL.scala 124:19]
    .io_in_0(m_626_io_in_0),
    .io_in_1(m_626_io_in_1),
    .io_out_0(m_626_io_out_0),
    .io_out_1(m_626_io_out_1)
  );
  Adder m_627 ( // @[MUL.scala 102:19]
    .io_x1(m_627_io_x1),
    .io_x2(m_627_io_x2),
    .io_x3(m_627_io_x3),
    .io_s(m_627_io_s),
    .io_cout(m_627_io_cout)
  );
  Adder m_628 ( // @[MUL.scala 102:19]
    .io_x1(m_628_io_x1),
    .io_x2(m_628_io_x2),
    .io_x3(m_628_io_x3),
    .io_s(m_628_io_s),
    .io_cout(m_628_io_cout)
  );
  Adder m_629 ( // @[MUL.scala 102:19]
    .io_x1(m_629_io_x1),
    .io_x2(m_629_io_x2),
    .io_x3(m_629_io_x3),
    .io_s(m_629_io_s),
    .io_cout(m_629_io_cout)
  );
  Adder m_630 ( // @[MUL.scala 102:19]
    .io_x1(m_630_io_x1),
    .io_x2(m_630_io_x2),
    .io_x3(m_630_io_x3),
    .io_s(m_630_io_s),
    .io_cout(m_630_io_cout)
  );
  Adder m_631 ( // @[MUL.scala 102:19]
    .io_x1(m_631_io_x1),
    .io_x2(m_631_io_x2),
    .io_x3(m_631_io_x3),
    .io_s(m_631_io_s),
    .io_cout(m_631_io_cout)
  );
  Adder m_632 ( // @[MUL.scala 102:19]
    .io_x1(m_632_io_x1),
    .io_x2(m_632_io_x2),
    .io_x3(m_632_io_x3),
    .io_s(m_632_io_s),
    .io_cout(m_632_io_cout)
  );
  Adder m_633 ( // @[MUL.scala 102:19]
    .io_x1(m_633_io_x1),
    .io_x2(m_633_io_x2),
    .io_x3(m_633_io_x3),
    .io_s(m_633_io_s),
    .io_cout(m_633_io_cout)
  );
  Half_Adder m_634 ( // @[MUL.scala 124:19]
    .io_in_0(m_634_io_in_0),
    .io_in_1(m_634_io_in_1),
    .io_out_0(m_634_io_out_0),
    .io_out_1(m_634_io_out_1)
  );
  Adder m_635 ( // @[MUL.scala 102:19]
    .io_x1(m_635_io_x1),
    .io_x2(m_635_io_x2),
    .io_x3(m_635_io_x3),
    .io_s(m_635_io_s),
    .io_cout(m_635_io_cout)
  );
  Adder m_636 ( // @[MUL.scala 102:19]
    .io_x1(m_636_io_x1),
    .io_x2(m_636_io_x2),
    .io_x3(m_636_io_x3),
    .io_s(m_636_io_s),
    .io_cout(m_636_io_cout)
  );
  Adder m_637 ( // @[MUL.scala 102:19]
    .io_x1(m_637_io_x1),
    .io_x2(m_637_io_x2),
    .io_x3(m_637_io_x3),
    .io_s(m_637_io_s),
    .io_cout(m_637_io_cout)
  );
  Adder m_638 ( // @[MUL.scala 102:19]
    .io_x1(m_638_io_x1),
    .io_x2(m_638_io_x2),
    .io_x3(m_638_io_x3),
    .io_s(m_638_io_s),
    .io_cout(m_638_io_cout)
  );
  Adder m_639 ( // @[MUL.scala 102:19]
    .io_x1(m_639_io_x1),
    .io_x2(m_639_io_x2),
    .io_x3(m_639_io_x3),
    .io_s(m_639_io_s),
    .io_cout(m_639_io_cout)
  );
  Adder m_640 ( // @[MUL.scala 102:19]
    .io_x1(m_640_io_x1),
    .io_x2(m_640_io_x2),
    .io_x3(m_640_io_x3),
    .io_s(m_640_io_s),
    .io_cout(m_640_io_cout)
  );
  Adder m_641 ( // @[MUL.scala 102:19]
    .io_x1(m_641_io_x1),
    .io_x2(m_641_io_x2),
    .io_x3(m_641_io_x3),
    .io_s(m_641_io_s),
    .io_cout(m_641_io_cout)
  );
  Adder m_642 ( // @[MUL.scala 102:19]
    .io_x1(m_642_io_x1),
    .io_x2(m_642_io_x2),
    .io_x3(m_642_io_x3),
    .io_s(m_642_io_s),
    .io_cout(m_642_io_cout)
  );
  Adder m_643 ( // @[MUL.scala 102:19]
    .io_x1(m_643_io_x1),
    .io_x2(m_643_io_x2),
    .io_x3(m_643_io_x3),
    .io_s(m_643_io_s),
    .io_cout(m_643_io_cout)
  );
  Adder m_644 ( // @[MUL.scala 102:19]
    .io_x1(m_644_io_x1),
    .io_x2(m_644_io_x2),
    .io_x3(m_644_io_x3),
    .io_s(m_644_io_s),
    .io_cout(m_644_io_cout)
  );
  Adder m_645 ( // @[MUL.scala 102:19]
    .io_x1(m_645_io_x1),
    .io_x2(m_645_io_x2),
    .io_x3(m_645_io_x3),
    .io_s(m_645_io_s),
    .io_cout(m_645_io_cout)
  );
  Adder m_646 ( // @[MUL.scala 102:19]
    .io_x1(m_646_io_x1),
    .io_x2(m_646_io_x2),
    .io_x3(m_646_io_x3),
    .io_s(m_646_io_s),
    .io_cout(m_646_io_cout)
  );
  Adder m_647 ( // @[MUL.scala 102:19]
    .io_x1(m_647_io_x1),
    .io_x2(m_647_io_x2),
    .io_x3(m_647_io_x3),
    .io_s(m_647_io_s),
    .io_cout(m_647_io_cout)
  );
  Adder m_648 ( // @[MUL.scala 102:19]
    .io_x1(m_648_io_x1),
    .io_x2(m_648_io_x2),
    .io_x3(m_648_io_x3),
    .io_s(m_648_io_s),
    .io_cout(m_648_io_cout)
  );
  Adder m_649 ( // @[MUL.scala 102:19]
    .io_x1(m_649_io_x1),
    .io_x2(m_649_io_x2),
    .io_x3(m_649_io_x3),
    .io_s(m_649_io_s),
    .io_cout(m_649_io_cout)
  );
  Adder m_650 ( // @[MUL.scala 102:19]
    .io_x1(m_650_io_x1),
    .io_x2(m_650_io_x2),
    .io_x3(m_650_io_x3),
    .io_s(m_650_io_s),
    .io_cout(m_650_io_cout)
  );
  Adder m_651 ( // @[MUL.scala 102:19]
    .io_x1(m_651_io_x1),
    .io_x2(m_651_io_x2),
    .io_x3(m_651_io_x3),
    .io_s(m_651_io_s),
    .io_cout(m_651_io_cout)
  );
  Adder m_652 ( // @[MUL.scala 102:19]
    .io_x1(m_652_io_x1),
    .io_x2(m_652_io_x2),
    .io_x3(m_652_io_x3),
    .io_s(m_652_io_s),
    .io_cout(m_652_io_cout)
  );
  Adder m_653 ( // @[MUL.scala 102:19]
    .io_x1(m_653_io_x1),
    .io_x2(m_653_io_x2),
    .io_x3(m_653_io_x3),
    .io_s(m_653_io_s),
    .io_cout(m_653_io_cout)
  );
  Adder m_654 ( // @[MUL.scala 102:19]
    .io_x1(m_654_io_x1),
    .io_x2(m_654_io_x2),
    .io_x3(m_654_io_x3),
    .io_s(m_654_io_s),
    .io_cout(m_654_io_cout)
  );
  Adder m_655 ( // @[MUL.scala 102:19]
    .io_x1(m_655_io_x1),
    .io_x2(m_655_io_x2),
    .io_x3(m_655_io_x3),
    .io_s(m_655_io_s),
    .io_cout(m_655_io_cout)
  );
  Adder m_656 ( // @[MUL.scala 102:19]
    .io_x1(m_656_io_x1),
    .io_x2(m_656_io_x2),
    .io_x3(m_656_io_x3),
    .io_s(m_656_io_s),
    .io_cout(m_656_io_cout)
  );
  Adder m_657 ( // @[MUL.scala 102:19]
    .io_x1(m_657_io_x1),
    .io_x2(m_657_io_x2),
    .io_x3(m_657_io_x3),
    .io_s(m_657_io_s),
    .io_cout(m_657_io_cout)
  );
  Adder m_658 ( // @[MUL.scala 102:19]
    .io_x1(m_658_io_x1),
    .io_x2(m_658_io_x2),
    .io_x3(m_658_io_x3),
    .io_s(m_658_io_s),
    .io_cout(m_658_io_cout)
  );
  Adder m_659 ( // @[MUL.scala 102:19]
    .io_x1(m_659_io_x1),
    .io_x2(m_659_io_x2),
    .io_x3(m_659_io_x3),
    .io_s(m_659_io_s),
    .io_cout(m_659_io_cout)
  );
  Adder m_660 ( // @[MUL.scala 102:19]
    .io_x1(m_660_io_x1),
    .io_x2(m_660_io_x2),
    .io_x3(m_660_io_x3),
    .io_s(m_660_io_s),
    .io_cout(m_660_io_cout)
  );
  Adder m_661 ( // @[MUL.scala 102:19]
    .io_x1(m_661_io_x1),
    .io_x2(m_661_io_x2),
    .io_x3(m_661_io_x3),
    .io_s(m_661_io_s),
    .io_cout(m_661_io_cout)
  );
  Adder m_662 ( // @[MUL.scala 102:19]
    .io_x1(m_662_io_x1),
    .io_x2(m_662_io_x2),
    .io_x3(m_662_io_x3),
    .io_s(m_662_io_s),
    .io_cout(m_662_io_cout)
  );
  Adder m_663 ( // @[MUL.scala 102:19]
    .io_x1(m_663_io_x1),
    .io_x2(m_663_io_x2),
    .io_x3(m_663_io_x3),
    .io_s(m_663_io_s),
    .io_cout(m_663_io_cout)
  );
  Adder m_664 ( // @[MUL.scala 102:19]
    .io_x1(m_664_io_x1),
    .io_x2(m_664_io_x2),
    .io_x3(m_664_io_x3),
    .io_s(m_664_io_s),
    .io_cout(m_664_io_cout)
  );
  Adder m_665 ( // @[MUL.scala 102:19]
    .io_x1(m_665_io_x1),
    .io_x2(m_665_io_x2),
    .io_x3(m_665_io_x3),
    .io_s(m_665_io_s),
    .io_cout(m_665_io_cout)
  );
  Adder m_666 ( // @[MUL.scala 102:19]
    .io_x1(m_666_io_x1),
    .io_x2(m_666_io_x2),
    .io_x3(m_666_io_x3),
    .io_s(m_666_io_s),
    .io_cout(m_666_io_cout)
  );
  Adder m_667 ( // @[MUL.scala 102:19]
    .io_x1(m_667_io_x1),
    .io_x2(m_667_io_x2),
    .io_x3(m_667_io_x3),
    .io_s(m_667_io_s),
    .io_cout(m_667_io_cout)
  );
  Adder m_668 ( // @[MUL.scala 102:19]
    .io_x1(m_668_io_x1),
    .io_x2(m_668_io_x2),
    .io_x3(m_668_io_x3),
    .io_s(m_668_io_s),
    .io_cout(m_668_io_cout)
  );
  Half_Adder m_669 ( // @[MUL.scala 124:19]
    .io_in_0(m_669_io_in_0),
    .io_in_1(m_669_io_in_1),
    .io_out_0(m_669_io_out_0),
    .io_out_1(m_669_io_out_1)
  );
  Adder m_670 ( // @[MUL.scala 102:19]
    .io_x1(m_670_io_x1),
    .io_x2(m_670_io_x2),
    .io_x3(m_670_io_x3),
    .io_s(m_670_io_s),
    .io_cout(m_670_io_cout)
  );
  Adder m_671 ( // @[MUL.scala 102:19]
    .io_x1(m_671_io_x1),
    .io_x2(m_671_io_x2),
    .io_x3(m_671_io_x3),
    .io_s(m_671_io_s),
    .io_cout(m_671_io_cout)
  );
  Adder m_672 ( // @[MUL.scala 102:19]
    .io_x1(m_672_io_x1),
    .io_x2(m_672_io_x2),
    .io_x3(m_672_io_x3),
    .io_s(m_672_io_s),
    .io_cout(m_672_io_cout)
  );
  Adder m_673 ( // @[MUL.scala 102:19]
    .io_x1(m_673_io_x1),
    .io_x2(m_673_io_x2),
    .io_x3(m_673_io_x3),
    .io_s(m_673_io_s),
    .io_cout(m_673_io_cout)
  );
  Adder m_674 ( // @[MUL.scala 102:19]
    .io_x1(m_674_io_x1),
    .io_x2(m_674_io_x2),
    .io_x3(m_674_io_x3),
    .io_s(m_674_io_s),
    .io_cout(m_674_io_cout)
  );
  Adder m_675 ( // @[MUL.scala 102:19]
    .io_x1(m_675_io_x1),
    .io_x2(m_675_io_x2),
    .io_x3(m_675_io_x3),
    .io_s(m_675_io_s),
    .io_cout(m_675_io_cout)
  );
  Half_Adder m_676 ( // @[MUL.scala 124:19]
    .io_in_0(m_676_io_in_0),
    .io_in_1(m_676_io_in_1),
    .io_out_0(m_676_io_out_0),
    .io_out_1(m_676_io_out_1)
  );
  Adder m_677 ( // @[MUL.scala 102:19]
    .io_x1(m_677_io_x1),
    .io_x2(m_677_io_x2),
    .io_x3(m_677_io_x3),
    .io_s(m_677_io_s),
    .io_cout(m_677_io_cout)
  );
  Adder m_678 ( // @[MUL.scala 102:19]
    .io_x1(m_678_io_x1),
    .io_x2(m_678_io_x2),
    .io_x3(m_678_io_x3),
    .io_s(m_678_io_s),
    .io_cout(m_678_io_cout)
  );
  Adder m_679 ( // @[MUL.scala 102:19]
    .io_x1(m_679_io_x1),
    .io_x2(m_679_io_x2),
    .io_x3(m_679_io_x3),
    .io_s(m_679_io_s),
    .io_cout(m_679_io_cout)
  );
  Adder m_680 ( // @[MUL.scala 102:19]
    .io_x1(m_680_io_x1),
    .io_x2(m_680_io_x2),
    .io_x3(m_680_io_x3),
    .io_s(m_680_io_s),
    .io_cout(m_680_io_cout)
  );
  Adder m_681 ( // @[MUL.scala 102:19]
    .io_x1(m_681_io_x1),
    .io_x2(m_681_io_x2),
    .io_x3(m_681_io_x3),
    .io_s(m_681_io_s),
    .io_cout(m_681_io_cout)
  );
  Adder m_682 ( // @[MUL.scala 102:19]
    .io_x1(m_682_io_x1),
    .io_x2(m_682_io_x2),
    .io_x3(m_682_io_x3),
    .io_s(m_682_io_s),
    .io_cout(m_682_io_cout)
  );
  Adder m_683 ( // @[MUL.scala 102:19]
    .io_x1(m_683_io_x1),
    .io_x2(m_683_io_x2),
    .io_x3(m_683_io_x3),
    .io_s(m_683_io_s),
    .io_cout(m_683_io_cout)
  );
  Adder m_684 ( // @[MUL.scala 102:19]
    .io_x1(m_684_io_x1),
    .io_x2(m_684_io_x2),
    .io_x3(m_684_io_x3),
    .io_s(m_684_io_s),
    .io_cout(m_684_io_cout)
  );
  Adder m_685 ( // @[MUL.scala 102:19]
    .io_x1(m_685_io_x1),
    .io_x2(m_685_io_x2),
    .io_x3(m_685_io_x3),
    .io_s(m_685_io_s),
    .io_cout(m_685_io_cout)
  );
  Adder m_686 ( // @[MUL.scala 102:19]
    .io_x1(m_686_io_x1),
    .io_x2(m_686_io_x2),
    .io_x3(m_686_io_x3),
    .io_s(m_686_io_s),
    .io_cout(m_686_io_cout)
  );
  Adder m_687 ( // @[MUL.scala 102:19]
    .io_x1(m_687_io_x1),
    .io_x2(m_687_io_x2),
    .io_x3(m_687_io_x3),
    .io_s(m_687_io_s),
    .io_cout(m_687_io_cout)
  );
  Adder m_688 ( // @[MUL.scala 102:19]
    .io_x1(m_688_io_x1),
    .io_x2(m_688_io_x2),
    .io_x3(m_688_io_x3),
    .io_s(m_688_io_s),
    .io_cout(m_688_io_cout)
  );
  Adder m_689 ( // @[MUL.scala 102:19]
    .io_x1(m_689_io_x1),
    .io_x2(m_689_io_x2),
    .io_x3(m_689_io_x3),
    .io_s(m_689_io_s),
    .io_cout(m_689_io_cout)
  );
  Adder m_690 ( // @[MUL.scala 102:19]
    .io_x1(m_690_io_x1),
    .io_x2(m_690_io_x2),
    .io_x3(m_690_io_x3),
    .io_s(m_690_io_s),
    .io_cout(m_690_io_cout)
  );
  Adder m_691 ( // @[MUL.scala 102:19]
    .io_x1(m_691_io_x1),
    .io_x2(m_691_io_x2),
    .io_x3(m_691_io_x3),
    .io_s(m_691_io_s),
    .io_cout(m_691_io_cout)
  );
  Adder m_692 ( // @[MUL.scala 102:19]
    .io_x1(m_692_io_x1),
    .io_x2(m_692_io_x2),
    .io_x3(m_692_io_x3),
    .io_s(m_692_io_s),
    .io_cout(m_692_io_cout)
  );
  Adder m_693 ( // @[MUL.scala 102:19]
    .io_x1(m_693_io_x1),
    .io_x2(m_693_io_x2),
    .io_x3(m_693_io_x3),
    .io_s(m_693_io_s),
    .io_cout(m_693_io_cout)
  );
  Adder m_694 ( // @[MUL.scala 102:19]
    .io_x1(m_694_io_x1),
    .io_x2(m_694_io_x2),
    .io_x3(m_694_io_x3),
    .io_s(m_694_io_s),
    .io_cout(m_694_io_cout)
  );
  Adder m_695 ( // @[MUL.scala 102:19]
    .io_x1(m_695_io_x1),
    .io_x2(m_695_io_x2),
    .io_x3(m_695_io_x3),
    .io_s(m_695_io_s),
    .io_cout(m_695_io_cout)
  );
  Adder m_696 ( // @[MUL.scala 102:19]
    .io_x1(m_696_io_x1),
    .io_x2(m_696_io_x2),
    .io_x3(m_696_io_x3),
    .io_s(m_696_io_s),
    .io_cout(m_696_io_cout)
  );
  Adder m_697 ( // @[MUL.scala 102:19]
    .io_x1(m_697_io_x1),
    .io_x2(m_697_io_x2),
    .io_x3(m_697_io_x3),
    .io_s(m_697_io_s),
    .io_cout(m_697_io_cout)
  );
  Adder m_698 ( // @[MUL.scala 102:19]
    .io_x1(m_698_io_x1),
    .io_x2(m_698_io_x2),
    .io_x3(m_698_io_x3),
    .io_s(m_698_io_s),
    .io_cout(m_698_io_cout)
  );
  Adder m_699 ( // @[MUL.scala 102:19]
    .io_x1(m_699_io_x1),
    .io_x2(m_699_io_x2),
    .io_x3(m_699_io_x3),
    .io_s(m_699_io_s),
    .io_cout(m_699_io_cout)
  );
  Adder m_700 ( // @[MUL.scala 102:19]
    .io_x1(m_700_io_x1),
    .io_x2(m_700_io_x2),
    .io_x3(m_700_io_x3),
    .io_s(m_700_io_s),
    .io_cout(m_700_io_cout)
  );
  Adder m_701 ( // @[MUL.scala 102:19]
    .io_x1(m_701_io_x1),
    .io_x2(m_701_io_x2),
    .io_x3(m_701_io_x3),
    .io_s(m_701_io_s),
    .io_cout(m_701_io_cout)
  );
  Adder m_702 ( // @[MUL.scala 102:19]
    .io_x1(m_702_io_x1),
    .io_x2(m_702_io_x2),
    .io_x3(m_702_io_x3),
    .io_s(m_702_io_s),
    .io_cout(m_702_io_cout)
  );
  Adder m_703 ( // @[MUL.scala 102:19]
    .io_x1(m_703_io_x1),
    .io_x2(m_703_io_x2),
    .io_x3(m_703_io_x3),
    .io_s(m_703_io_s),
    .io_cout(m_703_io_cout)
  );
  Adder m_704 ( // @[MUL.scala 102:19]
    .io_x1(m_704_io_x1),
    .io_x2(m_704_io_x2),
    .io_x3(m_704_io_x3),
    .io_s(m_704_io_s),
    .io_cout(m_704_io_cout)
  );
  Adder m_705 ( // @[MUL.scala 102:19]
    .io_x1(m_705_io_x1),
    .io_x2(m_705_io_x2),
    .io_x3(m_705_io_x3),
    .io_s(m_705_io_s),
    .io_cout(m_705_io_cout)
  );
  Half_Adder m_706 ( // @[MUL.scala 124:19]
    .io_in_0(m_706_io_in_0),
    .io_in_1(m_706_io_in_1),
    .io_out_0(m_706_io_out_0),
    .io_out_1(m_706_io_out_1)
  );
  Adder m_707 ( // @[MUL.scala 102:19]
    .io_x1(m_707_io_x1),
    .io_x2(m_707_io_x2),
    .io_x3(m_707_io_x3),
    .io_s(m_707_io_s),
    .io_cout(m_707_io_cout)
  );
  Adder m_708 ( // @[MUL.scala 102:19]
    .io_x1(m_708_io_x1),
    .io_x2(m_708_io_x2),
    .io_x3(m_708_io_x3),
    .io_s(m_708_io_s),
    .io_cout(m_708_io_cout)
  );
  Adder m_709 ( // @[MUL.scala 102:19]
    .io_x1(m_709_io_x1),
    .io_x2(m_709_io_x2),
    .io_x3(m_709_io_x3),
    .io_s(m_709_io_s),
    .io_cout(m_709_io_cout)
  );
  Adder m_710 ( // @[MUL.scala 102:19]
    .io_x1(m_710_io_x1),
    .io_x2(m_710_io_x2),
    .io_x3(m_710_io_x3),
    .io_s(m_710_io_s),
    .io_cout(m_710_io_cout)
  );
  Adder m_711 ( // @[MUL.scala 102:19]
    .io_x1(m_711_io_x1),
    .io_x2(m_711_io_x2),
    .io_x3(m_711_io_x3),
    .io_s(m_711_io_s),
    .io_cout(m_711_io_cout)
  );
  Half_Adder m_712 ( // @[MUL.scala 124:19]
    .io_in_0(m_712_io_in_0),
    .io_in_1(m_712_io_in_1),
    .io_out_0(m_712_io_out_0),
    .io_out_1(m_712_io_out_1)
  );
  Adder m_713 ( // @[MUL.scala 102:19]
    .io_x1(m_713_io_x1),
    .io_x2(m_713_io_x2),
    .io_x3(m_713_io_x3),
    .io_s(m_713_io_s),
    .io_cout(m_713_io_cout)
  );
  Adder m_714 ( // @[MUL.scala 102:19]
    .io_x1(m_714_io_x1),
    .io_x2(m_714_io_x2),
    .io_x3(m_714_io_x3),
    .io_s(m_714_io_s),
    .io_cout(m_714_io_cout)
  );
  Adder m_715 ( // @[MUL.scala 102:19]
    .io_x1(m_715_io_x1),
    .io_x2(m_715_io_x2),
    .io_x3(m_715_io_x3),
    .io_s(m_715_io_s),
    .io_cout(m_715_io_cout)
  );
  Adder m_716 ( // @[MUL.scala 102:19]
    .io_x1(m_716_io_x1),
    .io_x2(m_716_io_x2),
    .io_x3(m_716_io_x3),
    .io_s(m_716_io_s),
    .io_cout(m_716_io_cout)
  );
  Adder m_717 ( // @[MUL.scala 102:19]
    .io_x1(m_717_io_x1),
    .io_x2(m_717_io_x2),
    .io_x3(m_717_io_x3),
    .io_s(m_717_io_s),
    .io_cout(m_717_io_cout)
  );
  Adder m_718 ( // @[MUL.scala 102:19]
    .io_x1(m_718_io_x1),
    .io_x2(m_718_io_x2),
    .io_x3(m_718_io_x3),
    .io_s(m_718_io_s),
    .io_cout(m_718_io_cout)
  );
  Adder m_719 ( // @[MUL.scala 102:19]
    .io_x1(m_719_io_x1),
    .io_x2(m_719_io_x2),
    .io_x3(m_719_io_x3),
    .io_s(m_719_io_s),
    .io_cout(m_719_io_cout)
  );
  Adder m_720 ( // @[MUL.scala 102:19]
    .io_x1(m_720_io_x1),
    .io_x2(m_720_io_x2),
    .io_x3(m_720_io_x3),
    .io_s(m_720_io_s),
    .io_cout(m_720_io_cout)
  );
  Adder m_721 ( // @[MUL.scala 102:19]
    .io_x1(m_721_io_x1),
    .io_x2(m_721_io_x2),
    .io_x3(m_721_io_x3),
    .io_s(m_721_io_s),
    .io_cout(m_721_io_cout)
  );
  Adder m_722 ( // @[MUL.scala 102:19]
    .io_x1(m_722_io_x1),
    .io_x2(m_722_io_x2),
    .io_x3(m_722_io_x3),
    .io_s(m_722_io_s),
    .io_cout(m_722_io_cout)
  );
  Adder m_723 ( // @[MUL.scala 102:19]
    .io_x1(m_723_io_x1),
    .io_x2(m_723_io_x2),
    .io_x3(m_723_io_x3),
    .io_s(m_723_io_s),
    .io_cout(m_723_io_cout)
  );
  Adder m_724 ( // @[MUL.scala 102:19]
    .io_x1(m_724_io_x1),
    .io_x2(m_724_io_x2),
    .io_x3(m_724_io_x3),
    .io_s(m_724_io_s),
    .io_cout(m_724_io_cout)
  );
  Adder m_725 ( // @[MUL.scala 102:19]
    .io_x1(m_725_io_x1),
    .io_x2(m_725_io_x2),
    .io_x3(m_725_io_x3),
    .io_s(m_725_io_s),
    .io_cout(m_725_io_cout)
  );
  Adder m_726 ( // @[MUL.scala 102:19]
    .io_x1(m_726_io_x1),
    .io_x2(m_726_io_x2),
    .io_x3(m_726_io_x3),
    .io_s(m_726_io_s),
    .io_cout(m_726_io_cout)
  );
  Adder m_727 ( // @[MUL.scala 102:19]
    .io_x1(m_727_io_x1),
    .io_x2(m_727_io_x2),
    .io_x3(m_727_io_x3),
    .io_s(m_727_io_s),
    .io_cout(m_727_io_cout)
  );
  Adder m_728 ( // @[MUL.scala 102:19]
    .io_x1(m_728_io_x1),
    .io_x2(m_728_io_x2),
    .io_x3(m_728_io_x3),
    .io_s(m_728_io_s),
    .io_cout(m_728_io_cout)
  );
  Adder m_729 ( // @[MUL.scala 102:19]
    .io_x1(m_729_io_x1),
    .io_x2(m_729_io_x2),
    .io_x3(m_729_io_x3),
    .io_s(m_729_io_s),
    .io_cout(m_729_io_cout)
  );
  Adder m_730 ( // @[MUL.scala 102:19]
    .io_x1(m_730_io_x1),
    .io_x2(m_730_io_x2),
    .io_x3(m_730_io_x3),
    .io_s(m_730_io_s),
    .io_cout(m_730_io_cout)
  );
  Adder m_731 ( // @[MUL.scala 102:19]
    .io_x1(m_731_io_x1),
    .io_x2(m_731_io_x2),
    .io_x3(m_731_io_x3),
    .io_s(m_731_io_s),
    .io_cout(m_731_io_cout)
  );
  Adder m_732 ( // @[MUL.scala 102:19]
    .io_x1(m_732_io_x1),
    .io_x2(m_732_io_x2),
    .io_x3(m_732_io_x3),
    .io_s(m_732_io_s),
    .io_cout(m_732_io_cout)
  );
  Adder m_733 ( // @[MUL.scala 102:19]
    .io_x1(m_733_io_x1),
    .io_x2(m_733_io_x2),
    .io_x3(m_733_io_x3),
    .io_s(m_733_io_s),
    .io_cout(m_733_io_cout)
  );
  Adder m_734 ( // @[MUL.scala 102:19]
    .io_x1(m_734_io_x1),
    .io_x2(m_734_io_x2),
    .io_x3(m_734_io_x3),
    .io_s(m_734_io_s),
    .io_cout(m_734_io_cout)
  );
  Adder m_735 ( // @[MUL.scala 102:19]
    .io_x1(m_735_io_x1),
    .io_x2(m_735_io_x2),
    .io_x3(m_735_io_x3),
    .io_s(m_735_io_s),
    .io_cout(m_735_io_cout)
  );
  Adder m_736 ( // @[MUL.scala 102:19]
    .io_x1(m_736_io_x1),
    .io_x2(m_736_io_x2),
    .io_x3(m_736_io_x3),
    .io_s(m_736_io_s),
    .io_cout(m_736_io_cout)
  );
  Half_Adder m_737 ( // @[MUL.scala 124:19]
    .io_in_0(m_737_io_in_0),
    .io_in_1(m_737_io_in_1),
    .io_out_0(m_737_io_out_0),
    .io_out_1(m_737_io_out_1)
  );
  Adder m_738 ( // @[MUL.scala 102:19]
    .io_x1(m_738_io_x1),
    .io_x2(m_738_io_x2),
    .io_x3(m_738_io_x3),
    .io_s(m_738_io_s),
    .io_cout(m_738_io_cout)
  );
  Adder m_739 ( // @[MUL.scala 102:19]
    .io_x1(m_739_io_x1),
    .io_x2(m_739_io_x2),
    .io_x3(m_739_io_x3),
    .io_s(m_739_io_s),
    .io_cout(m_739_io_cout)
  );
  Adder m_740 ( // @[MUL.scala 102:19]
    .io_x1(m_740_io_x1),
    .io_x2(m_740_io_x2),
    .io_x3(m_740_io_x3),
    .io_s(m_740_io_s),
    .io_cout(m_740_io_cout)
  );
  Adder m_741 ( // @[MUL.scala 102:19]
    .io_x1(m_741_io_x1),
    .io_x2(m_741_io_x2),
    .io_x3(m_741_io_x3),
    .io_s(m_741_io_s),
    .io_cout(m_741_io_cout)
  );
  Half_Adder m_742 ( // @[MUL.scala 124:19]
    .io_in_0(m_742_io_in_0),
    .io_in_1(m_742_io_in_1),
    .io_out_0(m_742_io_out_0),
    .io_out_1(m_742_io_out_1)
  );
  Adder m_743 ( // @[MUL.scala 102:19]
    .io_x1(m_743_io_x1),
    .io_x2(m_743_io_x2),
    .io_x3(m_743_io_x3),
    .io_s(m_743_io_s),
    .io_cout(m_743_io_cout)
  );
  Adder m_744 ( // @[MUL.scala 102:19]
    .io_x1(m_744_io_x1),
    .io_x2(m_744_io_x2),
    .io_x3(m_744_io_x3),
    .io_s(m_744_io_s),
    .io_cout(m_744_io_cout)
  );
  Adder m_745 ( // @[MUL.scala 102:19]
    .io_x1(m_745_io_x1),
    .io_x2(m_745_io_x2),
    .io_x3(m_745_io_x3),
    .io_s(m_745_io_s),
    .io_cout(m_745_io_cout)
  );
  Adder m_746 ( // @[MUL.scala 102:19]
    .io_x1(m_746_io_x1),
    .io_x2(m_746_io_x2),
    .io_x3(m_746_io_x3),
    .io_s(m_746_io_s),
    .io_cout(m_746_io_cout)
  );
  Adder m_747 ( // @[MUL.scala 102:19]
    .io_x1(m_747_io_x1),
    .io_x2(m_747_io_x2),
    .io_x3(m_747_io_x3),
    .io_s(m_747_io_s),
    .io_cout(m_747_io_cout)
  );
  Adder m_748 ( // @[MUL.scala 102:19]
    .io_x1(m_748_io_x1),
    .io_x2(m_748_io_x2),
    .io_x3(m_748_io_x3),
    .io_s(m_748_io_s),
    .io_cout(m_748_io_cout)
  );
  Adder m_749 ( // @[MUL.scala 102:19]
    .io_x1(m_749_io_x1),
    .io_x2(m_749_io_x2),
    .io_x3(m_749_io_x3),
    .io_s(m_749_io_s),
    .io_cout(m_749_io_cout)
  );
  Adder m_750 ( // @[MUL.scala 102:19]
    .io_x1(m_750_io_x1),
    .io_x2(m_750_io_x2),
    .io_x3(m_750_io_x3),
    .io_s(m_750_io_s),
    .io_cout(m_750_io_cout)
  );
  Adder m_751 ( // @[MUL.scala 102:19]
    .io_x1(m_751_io_x1),
    .io_x2(m_751_io_x2),
    .io_x3(m_751_io_x3),
    .io_s(m_751_io_s),
    .io_cout(m_751_io_cout)
  );
  Adder m_752 ( // @[MUL.scala 102:19]
    .io_x1(m_752_io_x1),
    .io_x2(m_752_io_x2),
    .io_x3(m_752_io_x3),
    .io_s(m_752_io_s),
    .io_cout(m_752_io_cout)
  );
  Adder m_753 ( // @[MUL.scala 102:19]
    .io_x1(m_753_io_x1),
    .io_x2(m_753_io_x2),
    .io_x3(m_753_io_x3),
    .io_s(m_753_io_s),
    .io_cout(m_753_io_cout)
  );
  Adder m_754 ( // @[MUL.scala 102:19]
    .io_x1(m_754_io_x1),
    .io_x2(m_754_io_x2),
    .io_x3(m_754_io_x3),
    .io_s(m_754_io_s),
    .io_cout(m_754_io_cout)
  );
  Adder m_755 ( // @[MUL.scala 102:19]
    .io_x1(m_755_io_x1),
    .io_x2(m_755_io_x2),
    .io_x3(m_755_io_x3),
    .io_s(m_755_io_s),
    .io_cout(m_755_io_cout)
  );
  Adder m_756 ( // @[MUL.scala 102:19]
    .io_x1(m_756_io_x1),
    .io_x2(m_756_io_x2),
    .io_x3(m_756_io_x3),
    .io_s(m_756_io_s),
    .io_cout(m_756_io_cout)
  );
  Adder m_757 ( // @[MUL.scala 102:19]
    .io_x1(m_757_io_x1),
    .io_x2(m_757_io_x2),
    .io_x3(m_757_io_x3),
    .io_s(m_757_io_s),
    .io_cout(m_757_io_cout)
  );
  Adder m_758 ( // @[MUL.scala 102:19]
    .io_x1(m_758_io_x1),
    .io_x2(m_758_io_x2),
    .io_x3(m_758_io_x3),
    .io_s(m_758_io_s),
    .io_cout(m_758_io_cout)
  );
  Adder m_759 ( // @[MUL.scala 102:19]
    .io_x1(m_759_io_x1),
    .io_x2(m_759_io_x2),
    .io_x3(m_759_io_x3),
    .io_s(m_759_io_s),
    .io_cout(m_759_io_cout)
  );
  Adder m_760 ( // @[MUL.scala 102:19]
    .io_x1(m_760_io_x1),
    .io_x2(m_760_io_x2),
    .io_x3(m_760_io_x3),
    .io_s(m_760_io_s),
    .io_cout(m_760_io_cout)
  );
  Adder m_761 ( // @[MUL.scala 102:19]
    .io_x1(m_761_io_x1),
    .io_x2(m_761_io_x2),
    .io_x3(m_761_io_x3),
    .io_s(m_761_io_s),
    .io_cout(m_761_io_cout)
  );
  Half_Adder m_762 ( // @[MUL.scala 124:19]
    .io_in_0(m_762_io_in_0),
    .io_in_1(m_762_io_in_1),
    .io_out_0(m_762_io_out_0),
    .io_out_1(m_762_io_out_1)
  );
  Adder m_763 ( // @[MUL.scala 102:19]
    .io_x1(m_763_io_x1),
    .io_x2(m_763_io_x2),
    .io_x3(m_763_io_x3),
    .io_s(m_763_io_s),
    .io_cout(m_763_io_cout)
  );
  Adder m_764 ( // @[MUL.scala 102:19]
    .io_x1(m_764_io_x1),
    .io_x2(m_764_io_x2),
    .io_x3(m_764_io_x3),
    .io_s(m_764_io_s),
    .io_cout(m_764_io_cout)
  );
  Adder m_765 ( // @[MUL.scala 102:19]
    .io_x1(m_765_io_x1),
    .io_x2(m_765_io_x2),
    .io_x3(m_765_io_x3),
    .io_s(m_765_io_s),
    .io_cout(m_765_io_cout)
  );
  Half_Adder m_766 ( // @[MUL.scala 124:19]
    .io_in_0(m_766_io_in_0),
    .io_in_1(m_766_io_in_1),
    .io_out_0(m_766_io_out_0),
    .io_out_1(m_766_io_out_1)
  );
  Adder m_767 ( // @[MUL.scala 102:19]
    .io_x1(m_767_io_x1),
    .io_x2(m_767_io_x2),
    .io_x3(m_767_io_x3),
    .io_s(m_767_io_s),
    .io_cout(m_767_io_cout)
  );
  Adder m_768 ( // @[MUL.scala 102:19]
    .io_x1(m_768_io_x1),
    .io_x2(m_768_io_x2),
    .io_x3(m_768_io_x3),
    .io_s(m_768_io_s),
    .io_cout(m_768_io_cout)
  );
  Adder m_769 ( // @[MUL.scala 102:19]
    .io_x1(m_769_io_x1),
    .io_x2(m_769_io_x2),
    .io_x3(m_769_io_x3),
    .io_s(m_769_io_s),
    .io_cout(m_769_io_cout)
  );
  Adder m_770 ( // @[MUL.scala 102:19]
    .io_x1(m_770_io_x1),
    .io_x2(m_770_io_x2),
    .io_x3(m_770_io_x3),
    .io_s(m_770_io_s),
    .io_cout(m_770_io_cout)
  );
  Adder m_771 ( // @[MUL.scala 102:19]
    .io_x1(m_771_io_x1),
    .io_x2(m_771_io_x2),
    .io_x3(m_771_io_x3),
    .io_s(m_771_io_s),
    .io_cout(m_771_io_cout)
  );
  Adder m_772 ( // @[MUL.scala 102:19]
    .io_x1(m_772_io_x1),
    .io_x2(m_772_io_x2),
    .io_x3(m_772_io_x3),
    .io_s(m_772_io_s),
    .io_cout(m_772_io_cout)
  );
  Adder m_773 ( // @[MUL.scala 102:19]
    .io_x1(m_773_io_x1),
    .io_x2(m_773_io_x2),
    .io_x3(m_773_io_x3),
    .io_s(m_773_io_s),
    .io_cout(m_773_io_cout)
  );
  Adder m_774 ( // @[MUL.scala 102:19]
    .io_x1(m_774_io_x1),
    .io_x2(m_774_io_x2),
    .io_x3(m_774_io_x3),
    .io_s(m_774_io_s),
    .io_cout(m_774_io_cout)
  );
  Adder m_775 ( // @[MUL.scala 102:19]
    .io_x1(m_775_io_x1),
    .io_x2(m_775_io_x2),
    .io_x3(m_775_io_x3),
    .io_s(m_775_io_s),
    .io_cout(m_775_io_cout)
  );
  Adder m_776 ( // @[MUL.scala 102:19]
    .io_x1(m_776_io_x1),
    .io_x2(m_776_io_x2),
    .io_x3(m_776_io_x3),
    .io_s(m_776_io_s),
    .io_cout(m_776_io_cout)
  );
  Adder m_777 ( // @[MUL.scala 102:19]
    .io_x1(m_777_io_x1),
    .io_x2(m_777_io_x2),
    .io_x3(m_777_io_x3),
    .io_s(m_777_io_s),
    .io_cout(m_777_io_cout)
  );
  Adder m_778 ( // @[MUL.scala 102:19]
    .io_x1(m_778_io_x1),
    .io_x2(m_778_io_x2),
    .io_x3(m_778_io_x3),
    .io_s(m_778_io_s),
    .io_cout(m_778_io_cout)
  );
  Adder m_779 ( // @[MUL.scala 102:19]
    .io_x1(m_779_io_x1),
    .io_x2(m_779_io_x2),
    .io_x3(m_779_io_x3),
    .io_s(m_779_io_s),
    .io_cout(m_779_io_cout)
  );
  Adder m_780 ( // @[MUL.scala 102:19]
    .io_x1(m_780_io_x1),
    .io_x2(m_780_io_x2),
    .io_x3(m_780_io_x3),
    .io_s(m_780_io_s),
    .io_cout(m_780_io_cout)
  );
  Half_Adder m_781 ( // @[MUL.scala 124:19]
    .io_in_0(m_781_io_in_0),
    .io_in_1(m_781_io_in_1),
    .io_out_0(m_781_io_out_0),
    .io_out_1(m_781_io_out_1)
  );
  Adder m_782 ( // @[MUL.scala 102:19]
    .io_x1(m_782_io_x1),
    .io_x2(m_782_io_x2),
    .io_x3(m_782_io_x3),
    .io_s(m_782_io_s),
    .io_cout(m_782_io_cout)
  );
  Adder m_783 ( // @[MUL.scala 102:19]
    .io_x1(m_783_io_x1),
    .io_x2(m_783_io_x2),
    .io_x3(m_783_io_x3),
    .io_s(m_783_io_s),
    .io_cout(m_783_io_cout)
  );
  Half_Adder m_784 ( // @[MUL.scala 124:19]
    .io_in_0(m_784_io_in_0),
    .io_in_1(m_784_io_in_1),
    .io_out_0(m_784_io_out_0),
    .io_out_1(m_784_io_out_1)
  );
  Adder m_785 ( // @[MUL.scala 102:19]
    .io_x1(m_785_io_x1),
    .io_x2(m_785_io_x2),
    .io_x3(m_785_io_x3),
    .io_s(m_785_io_s),
    .io_cout(m_785_io_cout)
  );
  Adder m_786 ( // @[MUL.scala 102:19]
    .io_x1(m_786_io_x1),
    .io_x2(m_786_io_x2),
    .io_x3(m_786_io_x3),
    .io_s(m_786_io_s),
    .io_cout(m_786_io_cout)
  );
  Adder m_787 ( // @[MUL.scala 102:19]
    .io_x1(m_787_io_x1),
    .io_x2(m_787_io_x2),
    .io_x3(m_787_io_x3),
    .io_s(m_787_io_s),
    .io_cout(m_787_io_cout)
  );
  Adder m_788 ( // @[MUL.scala 102:19]
    .io_x1(m_788_io_x1),
    .io_x2(m_788_io_x2),
    .io_x3(m_788_io_x3),
    .io_s(m_788_io_s),
    .io_cout(m_788_io_cout)
  );
  Adder m_789 ( // @[MUL.scala 102:19]
    .io_x1(m_789_io_x1),
    .io_x2(m_789_io_x2),
    .io_x3(m_789_io_x3),
    .io_s(m_789_io_s),
    .io_cout(m_789_io_cout)
  );
  Adder m_790 ( // @[MUL.scala 102:19]
    .io_x1(m_790_io_x1),
    .io_x2(m_790_io_x2),
    .io_x3(m_790_io_x3),
    .io_s(m_790_io_s),
    .io_cout(m_790_io_cout)
  );
  Adder m_791 ( // @[MUL.scala 102:19]
    .io_x1(m_791_io_x1),
    .io_x2(m_791_io_x2),
    .io_x3(m_791_io_x3),
    .io_s(m_791_io_s),
    .io_cout(m_791_io_cout)
  );
  Adder m_792 ( // @[MUL.scala 102:19]
    .io_x1(m_792_io_x1),
    .io_x2(m_792_io_x2),
    .io_x3(m_792_io_x3),
    .io_s(m_792_io_s),
    .io_cout(m_792_io_cout)
  );
  Adder m_793 ( // @[MUL.scala 102:19]
    .io_x1(m_793_io_x1),
    .io_x2(m_793_io_x2),
    .io_x3(m_793_io_x3),
    .io_s(m_793_io_s),
    .io_cout(m_793_io_cout)
  );
  Half_Adder m_794 ( // @[MUL.scala 124:19]
    .io_in_0(m_794_io_in_0),
    .io_in_1(m_794_io_in_1),
    .io_out_0(m_794_io_out_0),
    .io_out_1(m_794_io_out_1)
  );
  Adder m_795 ( // @[MUL.scala 102:19]
    .io_x1(m_795_io_x1),
    .io_x2(m_795_io_x2),
    .io_x3(m_795_io_x3),
    .io_s(m_795_io_s),
    .io_cout(m_795_io_cout)
  );
  Half_Adder m_796 ( // @[MUL.scala 124:19]
    .io_in_0(m_796_io_in_0),
    .io_in_1(m_796_io_in_1),
    .io_out_0(m_796_io_out_0),
    .io_out_1(m_796_io_out_1)
  );
  Adder m_797 ( // @[MUL.scala 102:19]
    .io_x1(m_797_io_x1),
    .io_x2(m_797_io_x2),
    .io_x3(m_797_io_x3),
    .io_s(m_797_io_s),
    .io_cout(m_797_io_cout)
  );
  Adder m_798 ( // @[MUL.scala 102:19]
    .io_x1(m_798_io_x1),
    .io_x2(m_798_io_x2),
    .io_x3(m_798_io_x3),
    .io_s(m_798_io_s),
    .io_cout(m_798_io_cout)
  );
  Adder m_799 ( // @[MUL.scala 102:19]
    .io_x1(m_799_io_x1),
    .io_x2(m_799_io_x2),
    .io_x3(m_799_io_x3),
    .io_s(m_799_io_s),
    .io_cout(m_799_io_cout)
  );
  Adder m_800 ( // @[MUL.scala 102:19]
    .io_x1(m_800_io_x1),
    .io_x2(m_800_io_x2),
    .io_x3(m_800_io_x3),
    .io_s(m_800_io_s),
    .io_cout(m_800_io_cout)
  );
  Half_Adder m_801 ( // @[MUL.scala 124:19]
    .io_in_0(m_801_io_in_0),
    .io_in_1(m_801_io_in_1),
    .io_out_0(m_801_io_out_0),
    .io_out_1(m_801_io_out_1)
  );
  Half_Adder m_802 ( // @[MUL.scala 124:19]
    .io_in_0(m_802_io_in_0),
    .io_in_1(m_802_io_in_1),
    .io_out_0(m_802_io_out_0),
    .io_out_1(m_802_io_out_1)
  );
  Half_Adder m_803 ( // @[MUL.scala 124:19]
    .io_in_0(m_803_io_in_0),
    .io_in_1(m_803_io_in_1),
    .io_out_0(m_803_io_out_0),
    .io_out_1(m_803_io_out_1)
  );
  Half_Adder m_804 ( // @[MUL.scala 124:19]
    .io_in_0(m_804_io_in_0),
    .io_in_1(m_804_io_in_1),
    .io_out_0(m_804_io_out_0),
    .io_out_1(m_804_io_out_1)
  );
  Half_Adder m_805 ( // @[MUL.scala 124:19]
    .io_in_0(m_805_io_in_0),
    .io_in_1(m_805_io_in_1),
    .io_out_0(m_805_io_out_0),
    .io_out_1(m_805_io_out_1)
  );
  Adder m_806 ( // @[MUL.scala 102:19]
    .io_x1(m_806_io_x1),
    .io_x2(m_806_io_x2),
    .io_x3(m_806_io_x3),
    .io_s(m_806_io_s),
    .io_cout(m_806_io_cout)
  );
  Adder m_807 ( // @[MUL.scala 102:19]
    .io_x1(m_807_io_x1),
    .io_x2(m_807_io_x2),
    .io_x3(m_807_io_x3),
    .io_s(m_807_io_s),
    .io_cout(m_807_io_cout)
  );
  Adder m_808 ( // @[MUL.scala 102:19]
    .io_x1(m_808_io_x1),
    .io_x2(m_808_io_x2),
    .io_x3(m_808_io_x3),
    .io_s(m_808_io_s),
    .io_cout(m_808_io_cout)
  );
  Adder m_809 ( // @[MUL.scala 102:19]
    .io_x1(m_809_io_x1),
    .io_x2(m_809_io_x2),
    .io_x3(m_809_io_x3),
    .io_s(m_809_io_s),
    .io_cout(m_809_io_cout)
  );
  Adder m_810 ( // @[MUL.scala 102:19]
    .io_x1(m_810_io_x1),
    .io_x2(m_810_io_x2),
    .io_x3(m_810_io_x3),
    .io_s(m_810_io_s),
    .io_cout(m_810_io_cout)
  );
  Adder m_811 ( // @[MUL.scala 102:19]
    .io_x1(m_811_io_x1),
    .io_x2(m_811_io_x2),
    .io_x3(m_811_io_x3),
    .io_s(m_811_io_s),
    .io_cout(m_811_io_cout)
  );
  Adder m_812 ( // @[MUL.scala 102:19]
    .io_x1(m_812_io_x1),
    .io_x2(m_812_io_x2),
    .io_x3(m_812_io_x3),
    .io_s(m_812_io_s),
    .io_cout(m_812_io_cout)
  );
  Half_Adder m_813 ( // @[MUL.scala 124:19]
    .io_in_0(m_813_io_in_0),
    .io_in_1(m_813_io_in_1),
    .io_out_0(m_813_io_out_0),
    .io_out_1(m_813_io_out_1)
  );
  Adder m_814 ( // @[MUL.scala 102:19]
    .io_x1(m_814_io_x1),
    .io_x2(m_814_io_x2),
    .io_x3(m_814_io_x3),
    .io_s(m_814_io_s),
    .io_cout(m_814_io_cout)
  );
  Half_Adder m_815 ( // @[MUL.scala 124:19]
    .io_in_0(m_815_io_in_0),
    .io_in_1(m_815_io_in_1),
    .io_out_0(m_815_io_out_0),
    .io_out_1(m_815_io_out_1)
  );
  Adder m_816 ( // @[MUL.scala 102:19]
    .io_x1(m_816_io_x1),
    .io_x2(m_816_io_x2),
    .io_x3(m_816_io_x3),
    .io_s(m_816_io_s),
    .io_cout(m_816_io_cout)
  );
  Half_Adder m_817 ( // @[MUL.scala 124:19]
    .io_in_0(m_817_io_in_0),
    .io_in_1(m_817_io_in_1),
    .io_out_0(m_817_io_out_0),
    .io_out_1(m_817_io_out_1)
  );
  Adder m_818 ( // @[MUL.scala 102:19]
    .io_x1(m_818_io_x1),
    .io_x2(m_818_io_x2),
    .io_x3(m_818_io_x3),
    .io_s(m_818_io_s),
    .io_cout(m_818_io_cout)
  );
  Adder m_819 ( // @[MUL.scala 102:19]
    .io_x1(m_819_io_x1),
    .io_x2(m_819_io_x2),
    .io_x3(m_819_io_x3),
    .io_s(m_819_io_s),
    .io_cout(m_819_io_cout)
  );
  Adder m_820 ( // @[MUL.scala 102:19]
    .io_x1(m_820_io_x1),
    .io_x2(m_820_io_x2),
    .io_x3(m_820_io_x3),
    .io_s(m_820_io_s),
    .io_cout(m_820_io_cout)
  );
  Adder m_821 ( // @[MUL.scala 102:19]
    .io_x1(m_821_io_x1),
    .io_x2(m_821_io_x2),
    .io_x3(m_821_io_x3),
    .io_s(m_821_io_s),
    .io_cout(m_821_io_cout)
  );
  Adder m_822 ( // @[MUL.scala 102:19]
    .io_x1(m_822_io_x1),
    .io_x2(m_822_io_x2),
    .io_x3(m_822_io_x3),
    .io_s(m_822_io_s),
    .io_cout(m_822_io_cout)
  );
  Adder m_823 ( // @[MUL.scala 102:19]
    .io_x1(m_823_io_x1),
    .io_x2(m_823_io_x2),
    .io_x3(m_823_io_x3),
    .io_s(m_823_io_s),
    .io_cout(m_823_io_cout)
  );
  Adder m_824 ( // @[MUL.scala 102:19]
    .io_x1(m_824_io_x1),
    .io_x2(m_824_io_x2),
    .io_x3(m_824_io_x3),
    .io_s(m_824_io_s),
    .io_cout(m_824_io_cout)
  );
  Adder m_825 ( // @[MUL.scala 102:19]
    .io_x1(m_825_io_x1),
    .io_x2(m_825_io_x2),
    .io_x3(m_825_io_x3),
    .io_s(m_825_io_s),
    .io_cout(m_825_io_cout)
  );
  Adder m_826 ( // @[MUL.scala 102:19]
    .io_x1(m_826_io_x1),
    .io_x2(m_826_io_x2),
    .io_x3(m_826_io_x3),
    .io_s(m_826_io_s),
    .io_cout(m_826_io_cout)
  );
  Adder m_827 ( // @[MUL.scala 102:19]
    .io_x1(m_827_io_x1),
    .io_x2(m_827_io_x2),
    .io_x3(m_827_io_x3),
    .io_s(m_827_io_s),
    .io_cout(m_827_io_cout)
  );
  Adder m_828 ( // @[MUL.scala 102:19]
    .io_x1(m_828_io_x1),
    .io_x2(m_828_io_x2),
    .io_x3(m_828_io_x3),
    .io_s(m_828_io_s),
    .io_cout(m_828_io_cout)
  );
  Adder m_829 ( // @[MUL.scala 102:19]
    .io_x1(m_829_io_x1),
    .io_x2(m_829_io_x2),
    .io_x3(m_829_io_x3),
    .io_s(m_829_io_s),
    .io_cout(m_829_io_cout)
  );
  Adder m_830 ( // @[MUL.scala 102:19]
    .io_x1(m_830_io_x1),
    .io_x2(m_830_io_x2),
    .io_x3(m_830_io_x3),
    .io_s(m_830_io_s),
    .io_cout(m_830_io_cout)
  );
  Adder m_831 ( // @[MUL.scala 102:19]
    .io_x1(m_831_io_x1),
    .io_x2(m_831_io_x2),
    .io_x3(m_831_io_x3),
    .io_s(m_831_io_s),
    .io_cout(m_831_io_cout)
  );
  Half_Adder m_832 ( // @[MUL.scala 124:19]
    .io_in_0(m_832_io_in_0),
    .io_in_1(m_832_io_in_1),
    .io_out_0(m_832_io_out_0),
    .io_out_1(m_832_io_out_1)
  );
  Adder m_833 ( // @[MUL.scala 102:19]
    .io_x1(m_833_io_x1),
    .io_x2(m_833_io_x2),
    .io_x3(m_833_io_x3),
    .io_s(m_833_io_s),
    .io_cout(m_833_io_cout)
  );
  Adder m_834 ( // @[MUL.scala 102:19]
    .io_x1(m_834_io_x1),
    .io_x2(m_834_io_x2),
    .io_x3(m_834_io_x3),
    .io_s(m_834_io_s),
    .io_cout(m_834_io_cout)
  );
  Half_Adder m_835 ( // @[MUL.scala 124:19]
    .io_in_0(m_835_io_in_0),
    .io_in_1(m_835_io_in_1),
    .io_out_0(m_835_io_out_0),
    .io_out_1(m_835_io_out_1)
  );
  Adder m_836 ( // @[MUL.scala 102:19]
    .io_x1(m_836_io_x1),
    .io_x2(m_836_io_x2),
    .io_x3(m_836_io_x3),
    .io_s(m_836_io_s),
    .io_cout(m_836_io_cout)
  );
  Adder m_837 ( // @[MUL.scala 102:19]
    .io_x1(m_837_io_x1),
    .io_x2(m_837_io_x2),
    .io_x3(m_837_io_x3),
    .io_s(m_837_io_s),
    .io_cout(m_837_io_cout)
  );
  Half_Adder m_838 ( // @[MUL.scala 124:19]
    .io_in_0(m_838_io_in_0),
    .io_in_1(m_838_io_in_1),
    .io_out_0(m_838_io_out_0),
    .io_out_1(m_838_io_out_1)
  );
  Adder m_839 ( // @[MUL.scala 102:19]
    .io_x1(m_839_io_x1),
    .io_x2(m_839_io_x2),
    .io_x3(m_839_io_x3),
    .io_s(m_839_io_s),
    .io_cout(m_839_io_cout)
  );
  Adder m_840 ( // @[MUL.scala 102:19]
    .io_x1(m_840_io_x1),
    .io_x2(m_840_io_x2),
    .io_x3(m_840_io_x3),
    .io_s(m_840_io_s),
    .io_cout(m_840_io_cout)
  );
  Adder m_841 ( // @[MUL.scala 102:19]
    .io_x1(m_841_io_x1),
    .io_x2(m_841_io_x2),
    .io_x3(m_841_io_x3),
    .io_s(m_841_io_s),
    .io_cout(m_841_io_cout)
  );
  Adder m_842 ( // @[MUL.scala 102:19]
    .io_x1(m_842_io_x1),
    .io_x2(m_842_io_x2),
    .io_x3(m_842_io_x3),
    .io_s(m_842_io_s),
    .io_cout(m_842_io_cout)
  );
  Adder m_843 ( // @[MUL.scala 102:19]
    .io_x1(m_843_io_x1),
    .io_x2(m_843_io_x2),
    .io_x3(m_843_io_x3),
    .io_s(m_843_io_s),
    .io_cout(m_843_io_cout)
  );
  Adder m_844 ( // @[MUL.scala 102:19]
    .io_x1(m_844_io_x1),
    .io_x2(m_844_io_x2),
    .io_x3(m_844_io_x3),
    .io_s(m_844_io_s),
    .io_cout(m_844_io_cout)
  );
  Adder m_845 ( // @[MUL.scala 102:19]
    .io_x1(m_845_io_x1),
    .io_x2(m_845_io_x2),
    .io_x3(m_845_io_x3),
    .io_s(m_845_io_s),
    .io_cout(m_845_io_cout)
  );
  Adder m_846 ( // @[MUL.scala 102:19]
    .io_x1(m_846_io_x1),
    .io_x2(m_846_io_x2),
    .io_x3(m_846_io_x3),
    .io_s(m_846_io_s),
    .io_cout(m_846_io_cout)
  );
  Adder m_847 ( // @[MUL.scala 102:19]
    .io_x1(m_847_io_x1),
    .io_x2(m_847_io_x2),
    .io_x3(m_847_io_x3),
    .io_s(m_847_io_s),
    .io_cout(m_847_io_cout)
  );
  Adder m_848 ( // @[MUL.scala 102:19]
    .io_x1(m_848_io_x1),
    .io_x2(m_848_io_x2),
    .io_x3(m_848_io_x3),
    .io_s(m_848_io_s),
    .io_cout(m_848_io_cout)
  );
  Adder m_849 ( // @[MUL.scala 102:19]
    .io_x1(m_849_io_x1),
    .io_x2(m_849_io_x2),
    .io_x3(m_849_io_x3),
    .io_s(m_849_io_s),
    .io_cout(m_849_io_cout)
  );
  Adder m_850 ( // @[MUL.scala 102:19]
    .io_x1(m_850_io_x1),
    .io_x2(m_850_io_x2),
    .io_x3(m_850_io_x3),
    .io_s(m_850_io_s),
    .io_cout(m_850_io_cout)
  );
  Adder m_851 ( // @[MUL.scala 102:19]
    .io_x1(m_851_io_x1),
    .io_x2(m_851_io_x2),
    .io_x3(m_851_io_x3),
    .io_s(m_851_io_s),
    .io_cout(m_851_io_cout)
  );
  Adder m_852 ( // @[MUL.scala 102:19]
    .io_x1(m_852_io_x1),
    .io_x2(m_852_io_x2),
    .io_x3(m_852_io_x3),
    .io_s(m_852_io_s),
    .io_cout(m_852_io_cout)
  );
  Adder m_853 ( // @[MUL.scala 102:19]
    .io_x1(m_853_io_x1),
    .io_x2(m_853_io_x2),
    .io_x3(m_853_io_x3),
    .io_s(m_853_io_s),
    .io_cout(m_853_io_cout)
  );
  Adder m_854 ( // @[MUL.scala 102:19]
    .io_x1(m_854_io_x1),
    .io_x2(m_854_io_x2),
    .io_x3(m_854_io_x3),
    .io_s(m_854_io_s),
    .io_cout(m_854_io_cout)
  );
  Adder m_855 ( // @[MUL.scala 102:19]
    .io_x1(m_855_io_x1),
    .io_x2(m_855_io_x2),
    .io_x3(m_855_io_x3),
    .io_s(m_855_io_s),
    .io_cout(m_855_io_cout)
  );
  Adder m_856 ( // @[MUL.scala 102:19]
    .io_x1(m_856_io_x1),
    .io_x2(m_856_io_x2),
    .io_x3(m_856_io_x3),
    .io_s(m_856_io_s),
    .io_cout(m_856_io_cout)
  );
  Adder m_857 ( // @[MUL.scala 102:19]
    .io_x1(m_857_io_x1),
    .io_x2(m_857_io_x2),
    .io_x3(m_857_io_x3),
    .io_s(m_857_io_s),
    .io_cout(m_857_io_cout)
  );
  Adder m_858 ( // @[MUL.scala 102:19]
    .io_x1(m_858_io_x1),
    .io_x2(m_858_io_x2),
    .io_x3(m_858_io_x3),
    .io_s(m_858_io_s),
    .io_cout(m_858_io_cout)
  );
  Adder m_859 ( // @[MUL.scala 102:19]
    .io_x1(m_859_io_x1),
    .io_x2(m_859_io_x2),
    .io_x3(m_859_io_x3),
    .io_s(m_859_io_s),
    .io_cout(m_859_io_cout)
  );
  Half_Adder m_860 ( // @[MUL.scala 124:19]
    .io_in_0(m_860_io_in_0),
    .io_in_1(m_860_io_in_1),
    .io_out_0(m_860_io_out_0),
    .io_out_1(m_860_io_out_1)
  );
  Adder m_861 ( // @[MUL.scala 102:19]
    .io_x1(m_861_io_x1),
    .io_x2(m_861_io_x2),
    .io_x3(m_861_io_x3),
    .io_s(m_861_io_s),
    .io_cout(m_861_io_cout)
  );
  Adder m_862 ( // @[MUL.scala 102:19]
    .io_x1(m_862_io_x1),
    .io_x2(m_862_io_x2),
    .io_x3(m_862_io_x3),
    .io_s(m_862_io_s),
    .io_cout(m_862_io_cout)
  );
  Adder m_863 ( // @[MUL.scala 102:19]
    .io_x1(m_863_io_x1),
    .io_x2(m_863_io_x2),
    .io_x3(m_863_io_x3),
    .io_s(m_863_io_s),
    .io_cout(m_863_io_cout)
  );
  Half_Adder m_864 ( // @[MUL.scala 124:19]
    .io_in_0(m_864_io_in_0),
    .io_in_1(m_864_io_in_1),
    .io_out_0(m_864_io_out_0),
    .io_out_1(m_864_io_out_1)
  );
  Adder m_865 ( // @[MUL.scala 102:19]
    .io_x1(m_865_io_x1),
    .io_x2(m_865_io_x2),
    .io_x3(m_865_io_x3),
    .io_s(m_865_io_s),
    .io_cout(m_865_io_cout)
  );
  Adder m_866 ( // @[MUL.scala 102:19]
    .io_x1(m_866_io_x1),
    .io_x2(m_866_io_x2),
    .io_x3(m_866_io_x3),
    .io_s(m_866_io_s),
    .io_cout(m_866_io_cout)
  );
  Adder m_867 ( // @[MUL.scala 102:19]
    .io_x1(m_867_io_x1),
    .io_x2(m_867_io_x2),
    .io_x3(m_867_io_x3),
    .io_s(m_867_io_s),
    .io_cout(m_867_io_cout)
  );
  Half_Adder m_868 ( // @[MUL.scala 124:19]
    .io_in_0(m_868_io_in_0),
    .io_in_1(m_868_io_in_1),
    .io_out_0(m_868_io_out_0),
    .io_out_1(m_868_io_out_1)
  );
  Adder m_869 ( // @[MUL.scala 102:19]
    .io_x1(m_869_io_x1),
    .io_x2(m_869_io_x2),
    .io_x3(m_869_io_x3),
    .io_s(m_869_io_s),
    .io_cout(m_869_io_cout)
  );
  Adder m_870 ( // @[MUL.scala 102:19]
    .io_x1(m_870_io_x1),
    .io_x2(m_870_io_x2),
    .io_x3(m_870_io_x3),
    .io_s(m_870_io_s),
    .io_cout(m_870_io_cout)
  );
  Adder m_871 ( // @[MUL.scala 102:19]
    .io_x1(m_871_io_x1),
    .io_x2(m_871_io_x2),
    .io_x3(m_871_io_x3),
    .io_s(m_871_io_s),
    .io_cout(m_871_io_cout)
  );
  Adder m_872 ( // @[MUL.scala 102:19]
    .io_x1(m_872_io_x1),
    .io_x2(m_872_io_x2),
    .io_x3(m_872_io_x3),
    .io_s(m_872_io_s),
    .io_cout(m_872_io_cout)
  );
  Adder m_873 ( // @[MUL.scala 102:19]
    .io_x1(m_873_io_x1),
    .io_x2(m_873_io_x2),
    .io_x3(m_873_io_x3),
    .io_s(m_873_io_s),
    .io_cout(m_873_io_cout)
  );
  Adder m_874 ( // @[MUL.scala 102:19]
    .io_x1(m_874_io_x1),
    .io_x2(m_874_io_x2),
    .io_x3(m_874_io_x3),
    .io_s(m_874_io_s),
    .io_cout(m_874_io_cout)
  );
  Adder m_875 ( // @[MUL.scala 102:19]
    .io_x1(m_875_io_x1),
    .io_x2(m_875_io_x2),
    .io_x3(m_875_io_x3),
    .io_s(m_875_io_s),
    .io_cout(m_875_io_cout)
  );
  Adder m_876 ( // @[MUL.scala 102:19]
    .io_x1(m_876_io_x1),
    .io_x2(m_876_io_x2),
    .io_x3(m_876_io_x3),
    .io_s(m_876_io_s),
    .io_cout(m_876_io_cout)
  );
  Adder m_877 ( // @[MUL.scala 102:19]
    .io_x1(m_877_io_x1),
    .io_x2(m_877_io_x2),
    .io_x3(m_877_io_x3),
    .io_s(m_877_io_s),
    .io_cout(m_877_io_cout)
  );
  Adder m_878 ( // @[MUL.scala 102:19]
    .io_x1(m_878_io_x1),
    .io_x2(m_878_io_x2),
    .io_x3(m_878_io_x3),
    .io_s(m_878_io_s),
    .io_cout(m_878_io_cout)
  );
  Adder m_879 ( // @[MUL.scala 102:19]
    .io_x1(m_879_io_x1),
    .io_x2(m_879_io_x2),
    .io_x3(m_879_io_x3),
    .io_s(m_879_io_s),
    .io_cout(m_879_io_cout)
  );
  Adder m_880 ( // @[MUL.scala 102:19]
    .io_x1(m_880_io_x1),
    .io_x2(m_880_io_x2),
    .io_x3(m_880_io_x3),
    .io_s(m_880_io_s),
    .io_cout(m_880_io_cout)
  );
  Adder m_881 ( // @[MUL.scala 102:19]
    .io_x1(m_881_io_x1),
    .io_x2(m_881_io_x2),
    .io_x3(m_881_io_x3),
    .io_s(m_881_io_s),
    .io_cout(m_881_io_cout)
  );
  Adder m_882 ( // @[MUL.scala 102:19]
    .io_x1(m_882_io_x1),
    .io_x2(m_882_io_x2),
    .io_x3(m_882_io_x3),
    .io_s(m_882_io_s),
    .io_cout(m_882_io_cout)
  );
  Adder m_883 ( // @[MUL.scala 102:19]
    .io_x1(m_883_io_x1),
    .io_x2(m_883_io_x2),
    .io_x3(m_883_io_x3),
    .io_s(m_883_io_s),
    .io_cout(m_883_io_cout)
  );
  Adder m_884 ( // @[MUL.scala 102:19]
    .io_x1(m_884_io_x1),
    .io_x2(m_884_io_x2),
    .io_x3(m_884_io_x3),
    .io_s(m_884_io_s),
    .io_cout(m_884_io_cout)
  );
  Adder m_885 ( // @[MUL.scala 102:19]
    .io_x1(m_885_io_x1),
    .io_x2(m_885_io_x2),
    .io_x3(m_885_io_x3),
    .io_s(m_885_io_s),
    .io_cout(m_885_io_cout)
  );
  Adder m_886 ( // @[MUL.scala 102:19]
    .io_x1(m_886_io_x1),
    .io_x2(m_886_io_x2),
    .io_x3(m_886_io_x3),
    .io_s(m_886_io_s),
    .io_cout(m_886_io_cout)
  );
  Adder m_887 ( // @[MUL.scala 102:19]
    .io_x1(m_887_io_x1),
    .io_x2(m_887_io_x2),
    .io_x3(m_887_io_x3),
    .io_s(m_887_io_s),
    .io_cout(m_887_io_cout)
  );
  Adder m_888 ( // @[MUL.scala 102:19]
    .io_x1(m_888_io_x1),
    .io_x2(m_888_io_x2),
    .io_x3(m_888_io_x3),
    .io_s(m_888_io_s),
    .io_cout(m_888_io_cout)
  );
  Adder m_889 ( // @[MUL.scala 102:19]
    .io_x1(m_889_io_x1),
    .io_x2(m_889_io_x2),
    .io_x3(m_889_io_x3),
    .io_s(m_889_io_s),
    .io_cout(m_889_io_cout)
  );
  Adder m_890 ( // @[MUL.scala 102:19]
    .io_x1(m_890_io_x1),
    .io_x2(m_890_io_x2),
    .io_x3(m_890_io_x3),
    .io_s(m_890_io_s),
    .io_cout(m_890_io_cout)
  );
  Adder m_891 ( // @[MUL.scala 102:19]
    .io_x1(m_891_io_x1),
    .io_x2(m_891_io_x2),
    .io_x3(m_891_io_x3),
    .io_s(m_891_io_s),
    .io_cout(m_891_io_cout)
  );
  Adder m_892 ( // @[MUL.scala 102:19]
    .io_x1(m_892_io_x1),
    .io_x2(m_892_io_x2),
    .io_x3(m_892_io_x3),
    .io_s(m_892_io_s),
    .io_cout(m_892_io_cout)
  );
  Adder m_893 ( // @[MUL.scala 102:19]
    .io_x1(m_893_io_x1),
    .io_x2(m_893_io_x2),
    .io_x3(m_893_io_x3),
    .io_s(m_893_io_s),
    .io_cout(m_893_io_cout)
  );
  Adder m_894 ( // @[MUL.scala 102:19]
    .io_x1(m_894_io_x1),
    .io_x2(m_894_io_x2),
    .io_x3(m_894_io_x3),
    .io_s(m_894_io_s),
    .io_cout(m_894_io_cout)
  );
  Adder m_895 ( // @[MUL.scala 102:19]
    .io_x1(m_895_io_x1),
    .io_x2(m_895_io_x2),
    .io_x3(m_895_io_x3),
    .io_s(m_895_io_s),
    .io_cout(m_895_io_cout)
  );
  Adder m_896 ( // @[MUL.scala 102:19]
    .io_x1(m_896_io_x1),
    .io_x2(m_896_io_x2),
    .io_x3(m_896_io_x3),
    .io_s(m_896_io_s),
    .io_cout(m_896_io_cout)
  );
  Half_Adder m_897 ( // @[MUL.scala 124:19]
    .io_in_0(m_897_io_in_0),
    .io_in_1(m_897_io_in_1),
    .io_out_0(m_897_io_out_0),
    .io_out_1(m_897_io_out_1)
  );
  Adder m_898 ( // @[MUL.scala 102:19]
    .io_x1(m_898_io_x1),
    .io_x2(m_898_io_x2),
    .io_x3(m_898_io_x3),
    .io_s(m_898_io_s),
    .io_cout(m_898_io_cout)
  );
  Adder m_899 ( // @[MUL.scala 102:19]
    .io_x1(m_899_io_x1),
    .io_x2(m_899_io_x2),
    .io_x3(m_899_io_x3),
    .io_s(m_899_io_s),
    .io_cout(m_899_io_cout)
  );
  Adder m_900 ( // @[MUL.scala 102:19]
    .io_x1(m_900_io_x1),
    .io_x2(m_900_io_x2),
    .io_x3(m_900_io_x3),
    .io_s(m_900_io_s),
    .io_cout(m_900_io_cout)
  );
  Adder m_901 ( // @[MUL.scala 102:19]
    .io_x1(m_901_io_x1),
    .io_x2(m_901_io_x2),
    .io_x3(m_901_io_x3),
    .io_s(m_901_io_s),
    .io_cout(m_901_io_cout)
  );
  Half_Adder m_902 ( // @[MUL.scala 124:19]
    .io_in_0(m_902_io_in_0),
    .io_in_1(m_902_io_in_1),
    .io_out_0(m_902_io_out_0),
    .io_out_1(m_902_io_out_1)
  );
  Adder m_903 ( // @[MUL.scala 102:19]
    .io_x1(m_903_io_x1),
    .io_x2(m_903_io_x2),
    .io_x3(m_903_io_x3),
    .io_s(m_903_io_s),
    .io_cout(m_903_io_cout)
  );
  Adder m_904 ( // @[MUL.scala 102:19]
    .io_x1(m_904_io_x1),
    .io_x2(m_904_io_x2),
    .io_x3(m_904_io_x3),
    .io_s(m_904_io_s),
    .io_cout(m_904_io_cout)
  );
  Adder m_905 ( // @[MUL.scala 102:19]
    .io_x1(m_905_io_x1),
    .io_x2(m_905_io_x2),
    .io_x3(m_905_io_x3),
    .io_s(m_905_io_s),
    .io_cout(m_905_io_cout)
  );
  Adder m_906 ( // @[MUL.scala 102:19]
    .io_x1(m_906_io_x1),
    .io_x2(m_906_io_x2),
    .io_x3(m_906_io_x3),
    .io_s(m_906_io_s),
    .io_cout(m_906_io_cout)
  );
  Half_Adder m_907 ( // @[MUL.scala 124:19]
    .io_in_0(m_907_io_in_0),
    .io_in_1(m_907_io_in_1),
    .io_out_0(m_907_io_out_0),
    .io_out_1(m_907_io_out_1)
  );
  Adder m_908 ( // @[MUL.scala 102:19]
    .io_x1(m_908_io_x1),
    .io_x2(m_908_io_x2),
    .io_x3(m_908_io_x3),
    .io_s(m_908_io_s),
    .io_cout(m_908_io_cout)
  );
  Adder m_909 ( // @[MUL.scala 102:19]
    .io_x1(m_909_io_x1),
    .io_x2(m_909_io_x2),
    .io_x3(m_909_io_x3),
    .io_s(m_909_io_s),
    .io_cout(m_909_io_cout)
  );
  Adder m_910 ( // @[MUL.scala 102:19]
    .io_x1(m_910_io_x1),
    .io_x2(m_910_io_x2),
    .io_x3(m_910_io_x3),
    .io_s(m_910_io_s),
    .io_cout(m_910_io_cout)
  );
  Adder m_911 ( // @[MUL.scala 102:19]
    .io_x1(m_911_io_x1),
    .io_x2(m_911_io_x2),
    .io_x3(m_911_io_x3),
    .io_s(m_911_io_s),
    .io_cout(m_911_io_cout)
  );
  Adder m_912 ( // @[MUL.scala 102:19]
    .io_x1(m_912_io_x1),
    .io_x2(m_912_io_x2),
    .io_x3(m_912_io_x3),
    .io_s(m_912_io_s),
    .io_cout(m_912_io_cout)
  );
  Adder m_913 ( // @[MUL.scala 102:19]
    .io_x1(m_913_io_x1),
    .io_x2(m_913_io_x2),
    .io_x3(m_913_io_x3),
    .io_s(m_913_io_s),
    .io_cout(m_913_io_cout)
  );
  Adder m_914 ( // @[MUL.scala 102:19]
    .io_x1(m_914_io_x1),
    .io_x2(m_914_io_x2),
    .io_x3(m_914_io_x3),
    .io_s(m_914_io_s),
    .io_cout(m_914_io_cout)
  );
  Adder m_915 ( // @[MUL.scala 102:19]
    .io_x1(m_915_io_x1),
    .io_x2(m_915_io_x2),
    .io_x3(m_915_io_x3),
    .io_s(m_915_io_s),
    .io_cout(m_915_io_cout)
  );
  Adder m_916 ( // @[MUL.scala 102:19]
    .io_x1(m_916_io_x1),
    .io_x2(m_916_io_x2),
    .io_x3(m_916_io_x3),
    .io_s(m_916_io_s),
    .io_cout(m_916_io_cout)
  );
  Adder m_917 ( // @[MUL.scala 102:19]
    .io_x1(m_917_io_x1),
    .io_x2(m_917_io_x2),
    .io_x3(m_917_io_x3),
    .io_s(m_917_io_s),
    .io_cout(m_917_io_cout)
  );
  Adder m_918 ( // @[MUL.scala 102:19]
    .io_x1(m_918_io_x1),
    .io_x2(m_918_io_x2),
    .io_x3(m_918_io_x3),
    .io_s(m_918_io_s),
    .io_cout(m_918_io_cout)
  );
  Adder m_919 ( // @[MUL.scala 102:19]
    .io_x1(m_919_io_x1),
    .io_x2(m_919_io_x2),
    .io_x3(m_919_io_x3),
    .io_s(m_919_io_s),
    .io_cout(m_919_io_cout)
  );
  Adder m_920 ( // @[MUL.scala 102:19]
    .io_x1(m_920_io_x1),
    .io_x2(m_920_io_x2),
    .io_x3(m_920_io_x3),
    .io_s(m_920_io_s),
    .io_cout(m_920_io_cout)
  );
  Adder m_921 ( // @[MUL.scala 102:19]
    .io_x1(m_921_io_x1),
    .io_x2(m_921_io_x2),
    .io_x3(m_921_io_x3),
    .io_s(m_921_io_s),
    .io_cout(m_921_io_cout)
  );
  Adder m_922 ( // @[MUL.scala 102:19]
    .io_x1(m_922_io_x1),
    .io_x2(m_922_io_x2),
    .io_x3(m_922_io_x3),
    .io_s(m_922_io_s),
    .io_cout(m_922_io_cout)
  );
  Adder m_923 ( // @[MUL.scala 102:19]
    .io_x1(m_923_io_x1),
    .io_x2(m_923_io_x2),
    .io_x3(m_923_io_x3),
    .io_s(m_923_io_s),
    .io_cout(m_923_io_cout)
  );
  Adder m_924 ( // @[MUL.scala 102:19]
    .io_x1(m_924_io_x1),
    .io_x2(m_924_io_x2),
    .io_x3(m_924_io_x3),
    .io_s(m_924_io_s),
    .io_cout(m_924_io_cout)
  );
  Adder m_925 ( // @[MUL.scala 102:19]
    .io_x1(m_925_io_x1),
    .io_x2(m_925_io_x2),
    .io_x3(m_925_io_x3),
    .io_s(m_925_io_s),
    .io_cout(m_925_io_cout)
  );
  Adder m_926 ( // @[MUL.scala 102:19]
    .io_x1(m_926_io_x1),
    .io_x2(m_926_io_x2),
    .io_x3(m_926_io_x3),
    .io_s(m_926_io_s),
    .io_cout(m_926_io_cout)
  );
  Adder m_927 ( // @[MUL.scala 102:19]
    .io_x1(m_927_io_x1),
    .io_x2(m_927_io_x2),
    .io_x3(m_927_io_x3),
    .io_s(m_927_io_s),
    .io_cout(m_927_io_cout)
  );
  Adder m_928 ( // @[MUL.scala 102:19]
    .io_x1(m_928_io_x1),
    .io_x2(m_928_io_x2),
    .io_x3(m_928_io_x3),
    .io_s(m_928_io_s),
    .io_cout(m_928_io_cout)
  );
  Adder m_929 ( // @[MUL.scala 102:19]
    .io_x1(m_929_io_x1),
    .io_x2(m_929_io_x2),
    .io_x3(m_929_io_x3),
    .io_s(m_929_io_s),
    .io_cout(m_929_io_cout)
  );
  Adder m_930 ( // @[MUL.scala 102:19]
    .io_x1(m_930_io_x1),
    .io_x2(m_930_io_x2),
    .io_x3(m_930_io_x3),
    .io_s(m_930_io_s),
    .io_cout(m_930_io_cout)
  );
  Adder m_931 ( // @[MUL.scala 102:19]
    .io_x1(m_931_io_x1),
    .io_x2(m_931_io_x2),
    .io_x3(m_931_io_x3),
    .io_s(m_931_io_s),
    .io_cout(m_931_io_cout)
  );
  Adder m_932 ( // @[MUL.scala 102:19]
    .io_x1(m_932_io_x1),
    .io_x2(m_932_io_x2),
    .io_x3(m_932_io_x3),
    .io_s(m_932_io_s),
    .io_cout(m_932_io_cout)
  );
  Adder m_933 ( // @[MUL.scala 102:19]
    .io_x1(m_933_io_x1),
    .io_x2(m_933_io_x2),
    .io_x3(m_933_io_x3),
    .io_s(m_933_io_s),
    .io_cout(m_933_io_cout)
  );
  Adder m_934 ( // @[MUL.scala 102:19]
    .io_x1(m_934_io_x1),
    .io_x2(m_934_io_x2),
    .io_x3(m_934_io_x3),
    .io_s(m_934_io_s),
    .io_cout(m_934_io_cout)
  );
  Adder m_935 ( // @[MUL.scala 102:19]
    .io_x1(m_935_io_x1),
    .io_x2(m_935_io_x2),
    .io_x3(m_935_io_x3),
    .io_s(m_935_io_s),
    .io_cout(m_935_io_cout)
  );
  Adder m_936 ( // @[MUL.scala 102:19]
    .io_x1(m_936_io_x1),
    .io_x2(m_936_io_x2),
    .io_x3(m_936_io_x3),
    .io_s(m_936_io_s),
    .io_cout(m_936_io_cout)
  );
  Adder m_937 ( // @[MUL.scala 102:19]
    .io_x1(m_937_io_x1),
    .io_x2(m_937_io_x2),
    .io_x3(m_937_io_x3),
    .io_s(m_937_io_s),
    .io_cout(m_937_io_cout)
  );
  Adder m_938 ( // @[MUL.scala 102:19]
    .io_x1(m_938_io_x1),
    .io_x2(m_938_io_x2),
    .io_x3(m_938_io_x3),
    .io_s(m_938_io_s),
    .io_cout(m_938_io_cout)
  );
  Adder m_939 ( // @[MUL.scala 102:19]
    .io_x1(m_939_io_x1),
    .io_x2(m_939_io_x2),
    .io_x3(m_939_io_x3),
    .io_s(m_939_io_s),
    .io_cout(m_939_io_cout)
  );
  Adder m_940 ( // @[MUL.scala 102:19]
    .io_x1(m_940_io_x1),
    .io_x2(m_940_io_x2),
    .io_x3(m_940_io_x3),
    .io_s(m_940_io_s),
    .io_cout(m_940_io_cout)
  );
  Adder m_941 ( // @[MUL.scala 102:19]
    .io_x1(m_941_io_x1),
    .io_x2(m_941_io_x2),
    .io_x3(m_941_io_x3),
    .io_s(m_941_io_s),
    .io_cout(m_941_io_cout)
  );
  Adder m_942 ( // @[MUL.scala 102:19]
    .io_x1(m_942_io_x1),
    .io_x2(m_942_io_x2),
    .io_x3(m_942_io_x3),
    .io_s(m_942_io_s),
    .io_cout(m_942_io_cout)
  );
  Half_Adder m_943 ( // @[MUL.scala 124:19]
    .io_in_0(m_943_io_in_0),
    .io_in_1(m_943_io_in_1),
    .io_out_0(m_943_io_out_0),
    .io_out_1(m_943_io_out_1)
  );
  Adder m_944 ( // @[MUL.scala 102:19]
    .io_x1(m_944_io_x1),
    .io_x2(m_944_io_x2),
    .io_x3(m_944_io_x3),
    .io_s(m_944_io_s),
    .io_cout(m_944_io_cout)
  );
  Adder m_945 ( // @[MUL.scala 102:19]
    .io_x1(m_945_io_x1),
    .io_x2(m_945_io_x2),
    .io_x3(m_945_io_x3),
    .io_s(m_945_io_s),
    .io_cout(m_945_io_cout)
  );
  Adder m_946 ( // @[MUL.scala 102:19]
    .io_x1(m_946_io_x1),
    .io_x2(m_946_io_x2),
    .io_x3(m_946_io_x3),
    .io_s(m_946_io_s),
    .io_cout(m_946_io_cout)
  );
  Adder m_947 ( // @[MUL.scala 102:19]
    .io_x1(m_947_io_x1),
    .io_x2(m_947_io_x2),
    .io_x3(m_947_io_x3),
    .io_s(m_947_io_s),
    .io_cout(m_947_io_cout)
  );
  Adder m_948 ( // @[MUL.scala 102:19]
    .io_x1(m_948_io_x1),
    .io_x2(m_948_io_x2),
    .io_x3(m_948_io_x3),
    .io_s(m_948_io_s),
    .io_cout(m_948_io_cout)
  );
  Half_Adder m_949 ( // @[MUL.scala 124:19]
    .io_in_0(m_949_io_in_0),
    .io_in_1(m_949_io_in_1),
    .io_out_0(m_949_io_out_0),
    .io_out_1(m_949_io_out_1)
  );
  Adder m_950 ( // @[MUL.scala 102:19]
    .io_x1(m_950_io_x1),
    .io_x2(m_950_io_x2),
    .io_x3(m_950_io_x3),
    .io_s(m_950_io_s),
    .io_cout(m_950_io_cout)
  );
  Adder m_951 ( // @[MUL.scala 102:19]
    .io_x1(m_951_io_x1),
    .io_x2(m_951_io_x2),
    .io_x3(m_951_io_x3),
    .io_s(m_951_io_s),
    .io_cout(m_951_io_cout)
  );
  Adder m_952 ( // @[MUL.scala 102:19]
    .io_x1(m_952_io_x1),
    .io_x2(m_952_io_x2),
    .io_x3(m_952_io_x3),
    .io_s(m_952_io_s),
    .io_cout(m_952_io_cout)
  );
  Adder m_953 ( // @[MUL.scala 102:19]
    .io_x1(m_953_io_x1),
    .io_x2(m_953_io_x2),
    .io_x3(m_953_io_x3),
    .io_s(m_953_io_s),
    .io_cout(m_953_io_cout)
  );
  Adder m_954 ( // @[MUL.scala 102:19]
    .io_x1(m_954_io_x1),
    .io_x2(m_954_io_x2),
    .io_x3(m_954_io_x3),
    .io_s(m_954_io_s),
    .io_cout(m_954_io_cout)
  );
  Half_Adder m_955 ( // @[MUL.scala 124:19]
    .io_in_0(m_955_io_in_0),
    .io_in_1(m_955_io_in_1),
    .io_out_0(m_955_io_out_0),
    .io_out_1(m_955_io_out_1)
  );
  Adder m_956 ( // @[MUL.scala 102:19]
    .io_x1(m_956_io_x1),
    .io_x2(m_956_io_x2),
    .io_x3(m_956_io_x3),
    .io_s(m_956_io_s),
    .io_cout(m_956_io_cout)
  );
  Adder m_957 ( // @[MUL.scala 102:19]
    .io_x1(m_957_io_x1),
    .io_x2(m_957_io_x2),
    .io_x3(m_957_io_x3),
    .io_s(m_957_io_s),
    .io_cout(m_957_io_cout)
  );
  Adder m_958 ( // @[MUL.scala 102:19]
    .io_x1(m_958_io_x1),
    .io_x2(m_958_io_x2),
    .io_x3(m_958_io_x3),
    .io_s(m_958_io_s),
    .io_cout(m_958_io_cout)
  );
  Adder m_959 ( // @[MUL.scala 102:19]
    .io_x1(m_959_io_x1),
    .io_x2(m_959_io_x2),
    .io_x3(m_959_io_x3),
    .io_s(m_959_io_s),
    .io_cout(m_959_io_cout)
  );
  Adder m_960 ( // @[MUL.scala 102:19]
    .io_x1(m_960_io_x1),
    .io_x2(m_960_io_x2),
    .io_x3(m_960_io_x3),
    .io_s(m_960_io_s),
    .io_cout(m_960_io_cout)
  );
  Adder m_961 ( // @[MUL.scala 102:19]
    .io_x1(m_961_io_x1),
    .io_x2(m_961_io_x2),
    .io_x3(m_961_io_x3),
    .io_s(m_961_io_s),
    .io_cout(m_961_io_cout)
  );
  Adder m_962 ( // @[MUL.scala 102:19]
    .io_x1(m_962_io_x1),
    .io_x2(m_962_io_x2),
    .io_x3(m_962_io_x3),
    .io_s(m_962_io_s),
    .io_cout(m_962_io_cout)
  );
  Adder m_963 ( // @[MUL.scala 102:19]
    .io_x1(m_963_io_x1),
    .io_x2(m_963_io_x2),
    .io_x3(m_963_io_x3),
    .io_s(m_963_io_s),
    .io_cout(m_963_io_cout)
  );
  Adder m_964 ( // @[MUL.scala 102:19]
    .io_x1(m_964_io_x1),
    .io_x2(m_964_io_x2),
    .io_x3(m_964_io_x3),
    .io_s(m_964_io_s),
    .io_cout(m_964_io_cout)
  );
  Adder m_965 ( // @[MUL.scala 102:19]
    .io_x1(m_965_io_x1),
    .io_x2(m_965_io_x2),
    .io_x3(m_965_io_x3),
    .io_s(m_965_io_s),
    .io_cout(m_965_io_cout)
  );
  Adder m_966 ( // @[MUL.scala 102:19]
    .io_x1(m_966_io_x1),
    .io_x2(m_966_io_x2),
    .io_x3(m_966_io_x3),
    .io_s(m_966_io_s),
    .io_cout(m_966_io_cout)
  );
  Adder m_967 ( // @[MUL.scala 102:19]
    .io_x1(m_967_io_x1),
    .io_x2(m_967_io_x2),
    .io_x3(m_967_io_x3),
    .io_s(m_967_io_s),
    .io_cout(m_967_io_cout)
  );
  Adder m_968 ( // @[MUL.scala 102:19]
    .io_x1(m_968_io_x1),
    .io_x2(m_968_io_x2),
    .io_x3(m_968_io_x3),
    .io_s(m_968_io_s),
    .io_cout(m_968_io_cout)
  );
  Adder m_969 ( // @[MUL.scala 102:19]
    .io_x1(m_969_io_x1),
    .io_x2(m_969_io_x2),
    .io_x3(m_969_io_x3),
    .io_s(m_969_io_s),
    .io_cout(m_969_io_cout)
  );
  Adder m_970 ( // @[MUL.scala 102:19]
    .io_x1(m_970_io_x1),
    .io_x2(m_970_io_x2),
    .io_x3(m_970_io_x3),
    .io_s(m_970_io_s),
    .io_cout(m_970_io_cout)
  );
  Adder m_971 ( // @[MUL.scala 102:19]
    .io_x1(m_971_io_x1),
    .io_x2(m_971_io_x2),
    .io_x3(m_971_io_x3),
    .io_s(m_971_io_s),
    .io_cout(m_971_io_cout)
  );
  Adder m_972 ( // @[MUL.scala 102:19]
    .io_x1(m_972_io_x1),
    .io_x2(m_972_io_x2),
    .io_x3(m_972_io_x3),
    .io_s(m_972_io_s),
    .io_cout(m_972_io_cout)
  );
  Adder m_973 ( // @[MUL.scala 102:19]
    .io_x1(m_973_io_x1),
    .io_x2(m_973_io_x2),
    .io_x3(m_973_io_x3),
    .io_s(m_973_io_s),
    .io_cout(m_973_io_cout)
  );
  Adder m_974 ( // @[MUL.scala 102:19]
    .io_x1(m_974_io_x1),
    .io_x2(m_974_io_x2),
    .io_x3(m_974_io_x3),
    .io_s(m_974_io_s),
    .io_cout(m_974_io_cout)
  );
  Adder m_975 ( // @[MUL.scala 102:19]
    .io_x1(m_975_io_x1),
    .io_x2(m_975_io_x2),
    .io_x3(m_975_io_x3),
    .io_s(m_975_io_s),
    .io_cout(m_975_io_cout)
  );
  Adder m_976 ( // @[MUL.scala 102:19]
    .io_x1(m_976_io_x1),
    .io_x2(m_976_io_x2),
    .io_x3(m_976_io_x3),
    .io_s(m_976_io_s),
    .io_cout(m_976_io_cout)
  );
  Adder m_977 ( // @[MUL.scala 102:19]
    .io_x1(m_977_io_x1),
    .io_x2(m_977_io_x2),
    .io_x3(m_977_io_x3),
    .io_s(m_977_io_s),
    .io_cout(m_977_io_cout)
  );
  Adder m_978 ( // @[MUL.scala 102:19]
    .io_x1(m_978_io_x1),
    .io_x2(m_978_io_x2),
    .io_x3(m_978_io_x3),
    .io_s(m_978_io_s),
    .io_cout(m_978_io_cout)
  );
  Adder m_979 ( // @[MUL.scala 102:19]
    .io_x1(m_979_io_x1),
    .io_x2(m_979_io_x2),
    .io_x3(m_979_io_x3),
    .io_s(m_979_io_s),
    .io_cout(m_979_io_cout)
  );
  Adder m_980 ( // @[MUL.scala 102:19]
    .io_x1(m_980_io_x1),
    .io_x2(m_980_io_x2),
    .io_x3(m_980_io_x3),
    .io_s(m_980_io_s),
    .io_cout(m_980_io_cout)
  );
  Adder m_981 ( // @[MUL.scala 102:19]
    .io_x1(m_981_io_x1),
    .io_x2(m_981_io_x2),
    .io_x3(m_981_io_x3),
    .io_s(m_981_io_s),
    .io_cout(m_981_io_cout)
  );
  Adder m_982 ( // @[MUL.scala 102:19]
    .io_x1(m_982_io_x1),
    .io_x2(m_982_io_x2),
    .io_x3(m_982_io_x3),
    .io_s(m_982_io_s),
    .io_cout(m_982_io_cout)
  );
  Adder m_983 ( // @[MUL.scala 102:19]
    .io_x1(m_983_io_x1),
    .io_x2(m_983_io_x2),
    .io_x3(m_983_io_x3),
    .io_s(m_983_io_s),
    .io_cout(m_983_io_cout)
  );
  Adder m_984 ( // @[MUL.scala 102:19]
    .io_x1(m_984_io_x1),
    .io_x2(m_984_io_x2),
    .io_x3(m_984_io_x3),
    .io_s(m_984_io_s),
    .io_cout(m_984_io_cout)
  );
  Adder m_985 ( // @[MUL.scala 102:19]
    .io_x1(m_985_io_x1),
    .io_x2(m_985_io_x2),
    .io_x3(m_985_io_x3),
    .io_s(m_985_io_s),
    .io_cout(m_985_io_cout)
  );
  Adder m_986 ( // @[MUL.scala 102:19]
    .io_x1(m_986_io_x1),
    .io_x2(m_986_io_x2),
    .io_x3(m_986_io_x3),
    .io_s(m_986_io_s),
    .io_cout(m_986_io_cout)
  );
  Adder m_987 ( // @[MUL.scala 102:19]
    .io_x1(m_987_io_x1),
    .io_x2(m_987_io_x2),
    .io_x3(m_987_io_x3),
    .io_s(m_987_io_s),
    .io_cout(m_987_io_cout)
  );
  Adder m_988 ( // @[MUL.scala 102:19]
    .io_x1(m_988_io_x1),
    .io_x2(m_988_io_x2),
    .io_x3(m_988_io_x3),
    .io_s(m_988_io_s),
    .io_cout(m_988_io_cout)
  );
  Adder m_989 ( // @[MUL.scala 102:19]
    .io_x1(m_989_io_x1),
    .io_x2(m_989_io_x2),
    .io_x3(m_989_io_x3),
    .io_s(m_989_io_s),
    .io_cout(m_989_io_cout)
  );
  Adder m_990 ( // @[MUL.scala 102:19]
    .io_x1(m_990_io_x1),
    .io_x2(m_990_io_x2),
    .io_x3(m_990_io_x3),
    .io_s(m_990_io_s),
    .io_cout(m_990_io_cout)
  );
  Adder m_991 ( // @[MUL.scala 102:19]
    .io_x1(m_991_io_x1),
    .io_x2(m_991_io_x2),
    .io_x3(m_991_io_x3),
    .io_s(m_991_io_s),
    .io_cout(m_991_io_cout)
  );
  Adder m_992 ( // @[MUL.scala 102:19]
    .io_x1(m_992_io_x1),
    .io_x2(m_992_io_x2),
    .io_x3(m_992_io_x3),
    .io_s(m_992_io_s),
    .io_cout(m_992_io_cout)
  );
  Adder m_993 ( // @[MUL.scala 102:19]
    .io_x1(m_993_io_x1),
    .io_x2(m_993_io_x2),
    .io_x3(m_993_io_x3),
    .io_s(m_993_io_s),
    .io_cout(m_993_io_cout)
  );
  Adder m_994 ( // @[MUL.scala 102:19]
    .io_x1(m_994_io_x1),
    .io_x2(m_994_io_x2),
    .io_x3(m_994_io_x3),
    .io_s(m_994_io_s),
    .io_cout(m_994_io_cout)
  );
  Adder m_995 ( // @[MUL.scala 102:19]
    .io_x1(m_995_io_x1),
    .io_x2(m_995_io_x2),
    .io_x3(m_995_io_x3),
    .io_s(m_995_io_s),
    .io_cout(m_995_io_cout)
  );
  Adder m_996 ( // @[MUL.scala 102:19]
    .io_x1(m_996_io_x1),
    .io_x2(m_996_io_x2),
    .io_x3(m_996_io_x3),
    .io_s(m_996_io_s),
    .io_cout(m_996_io_cout)
  );
  Adder m_997 ( // @[MUL.scala 102:19]
    .io_x1(m_997_io_x1),
    .io_x2(m_997_io_x2),
    .io_x3(m_997_io_x3),
    .io_s(m_997_io_s),
    .io_cout(m_997_io_cout)
  );
  Half_Adder m_998 ( // @[MUL.scala 124:19]
    .io_in_0(m_998_io_in_0),
    .io_in_1(m_998_io_in_1),
    .io_out_0(m_998_io_out_0),
    .io_out_1(m_998_io_out_1)
  );
  Adder m_999 ( // @[MUL.scala 102:19]
    .io_x1(m_999_io_x1),
    .io_x2(m_999_io_x2),
    .io_x3(m_999_io_x3),
    .io_s(m_999_io_s),
    .io_cout(m_999_io_cout)
  );
  Adder m_1000 ( // @[MUL.scala 102:19]
    .io_x1(m_1000_io_x1),
    .io_x2(m_1000_io_x2),
    .io_x3(m_1000_io_x3),
    .io_s(m_1000_io_s),
    .io_cout(m_1000_io_cout)
  );
  Adder m_1001 ( // @[MUL.scala 102:19]
    .io_x1(m_1001_io_x1),
    .io_x2(m_1001_io_x2),
    .io_x3(m_1001_io_x3),
    .io_s(m_1001_io_s),
    .io_cout(m_1001_io_cout)
  );
  Adder m_1002 ( // @[MUL.scala 102:19]
    .io_x1(m_1002_io_x1),
    .io_x2(m_1002_io_x2),
    .io_x3(m_1002_io_x3),
    .io_s(m_1002_io_s),
    .io_cout(m_1002_io_cout)
  );
  Adder m_1003 ( // @[MUL.scala 102:19]
    .io_x1(m_1003_io_x1),
    .io_x2(m_1003_io_x2),
    .io_x3(m_1003_io_x3),
    .io_s(m_1003_io_s),
    .io_cout(m_1003_io_cout)
  );
  Adder m_1004 ( // @[MUL.scala 102:19]
    .io_x1(m_1004_io_x1),
    .io_x2(m_1004_io_x2),
    .io_x3(m_1004_io_x3),
    .io_s(m_1004_io_s),
    .io_cout(m_1004_io_cout)
  );
  Half_Adder m_1005 ( // @[MUL.scala 124:19]
    .io_in_0(m_1005_io_in_0),
    .io_in_1(m_1005_io_in_1),
    .io_out_0(m_1005_io_out_0),
    .io_out_1(m_1005_io_out_1)
  );
  Adder m_1006 ( // @[MUL.scala 102:19]
    .io_x1(m_1006_io_x1),
    .io_x2(m_1006_io_x2),
    .io_x3(m_1006_io_x3),
    .io_s(m_1006_io_s),
    .io_cout(m_1006_io_cout)
  );
  Adder m_1007 ( // @[MUL.scala 102:19]
    .io_x1(m_1007_io_x1),
    .io_x2(m_1007_io_x2),
    .io_x3(m_1007_io_x3),
    .io_s(m_1007_io_s),
    .io_cout(m_1007_io_cout)
  );
  Adder m_1008 ( // @[MUL.scala 102:19]
    .io_x1(m_1008_io_x1),
    .io_x2(m_1008_io_x2),
    .io_x3(m_1008_io_x3),
    .io_s(m_1008_io_s),
    .io_cout(m_1008_io_cout)
  );
  Adder m_1009 ( // @[MUL.scala 102:19]
    .io_x1(m_1009_io_x1),
    .io_x2(m_1009_io_x2),
    .io_x3(m_1009_io_x3),
    .io_s(m_1009_io_s),
    .io_cout(m_1009_io_cout)
  );
  Adder m_1010 ( // @[MUL.scala 102:19]
    .io_x1(m_1010_io_x1),
    .io_x2(m_1010_io_x2),
    .io_x3(m_1010_io_x3),
    .io_s(m_1010_io_s),
    .io_cout(m_1010_io_cout)
  );
  Adder m_1011 ( // @[MUL.scala 102:19]
    .io_x1(m_1011_io_x1),
    .io_x2(m_1011_io_x2),
    .io_x3(m_1011_io_x3),
    .io_s(m_1011_io_s),
    .io_cout(m_1011_io_cout)
  );
  Half_Adder m_1012 ( // @[MUL.scala 124:19]
    .io_in_0(m_1012_io_in_0),
    .io_in_1(m_1012_io_in_1),
    .io_out_0(m_1012_io_out_0),
    .io_out_1(m_1012_io_out_1)
  );
  Adder m_1013 ( // @[MUL.scala 102:19]
    .io_x1(m_1013_io_x1),
    .io_x2(m_1013_io_x2),
    .io_x3(m_1013_io_x3),
    .io_s(m_1013_io_s),
    .io_cout(m_1013_io_cout)
  );
  Adder m_1014 ( // @[MUL.scala 102:19]
    .io_x1(m_1014_io_x1),
    .io_x2(m_1014_io_x2),
    .io_x3(m_1014_io_x3),
    .io_s(m_1014_io_s),
    .io_cout(m_1014_io_cout)
  );
  Adder m_1015 ( // @[MUL.scala 102:19]
    .io_x1(m_1015_io_x1),
    .io_x2(m_1015_io_x2),
    .io_x3(m_1015_io_x3),
    .io_s(m_1015_io_s),
    .io_cout(m_1015_io_cout)
  );
  Adder m_1016 ( // @[MUL.scala 102:19]
    .io_x1(m_1016_io_x1),
    .io_x2(m_1016_io_x2),
    .io_x3(m_1016_io_x3),
    .io_s(m_1016_io_s),
    .io_cout(m_1016_io_cout)
  );
  Adder m_1017 ( // @[MUL.scala 102:19]
    .io_x1(m_1017_io_x1),
    .io_x2(m_1017_io_x2),
    .io_x3(m_1017_io_x3),
    .io_s(m_1017_io_s),
    .io_cout(m_1017_io_cout)
  );
  Adder m_1018 ( // @[MUL.scala 102:19]
    .io_x1(m_1018_io_x1),
    .io_x2(m_1018_io_x2),
    .io_x3(m_1018_io_x3),
    .io_s(m_1018_io_s),
    .io_cout(m_1018_io_cout)
  );
  Adder m_1019 ( // @[MUL.scala 102:19]
    .io_x1(m_1019_io_x1),
    .io_x2(m_1019_io_x2),
    .io_x3(m_1019_io_x3),
    .io_s(m_1019_io_s),
    .io_cout(m_1019_io_cout)
  );
  Adder m_1020 ( // @[MUL.scala 102:19]
    .io_x1(m_1020_io_x1),
    .io_x2(m_1020_io_x2),
    .io_x3(m_1020_io_x3),
    .io_s(m_1020_io_s),
    .io_cout(m_1020_io_cout)
  );
  Adder m_1021 ( // @[MUL.scala 102:19]
    .io_x1(m_1021_io_x1),
    .io_x2(m_1021_io_x2),
    .io_x3(m_1021_io_x3),
    .io_s(m_1021_io_s),
    .io_cout(m_1021_io_cout)
  );
  Adder m_1022 ( // @[MUL.scala 102:19]
    .io_x1(m_1022_io_x1),
    .io_x2(m_1022_io_x2),
    .io_x3(m_1022_io_x3),
    .io_s(m_1022_io_s),
    .io_cout(m_1022_io_cout)
  );
  Adder m_1023 ( // @[MUL.scala 102:19]
    .io_x1(m_1023_io_x1),
    .io_x2(m_1023_io_x2),
    .io_x3(m_1023_io_x3),
    .io_s(m_1023_io_s),
    .io_cout(m_1023_io_cout)
  );
  Adder m_1024 ( // @[MUL.scala 102:19]
    .io_x1(m_1024_io_x1),
    .io_x2(m_1024_io_x2),
    .io_x3(m_1024_io_x3),
    .io_s(m_1024_io_s),
    .io_cout(m_1024_io_cout)
  );
  Adder m_1025 ( // @[MUL.scala 102:19]
    .io_x1(m_1025_io_x1),
    .io_x2(m_1025_io_x2),
    .io_x3(m_1025_io_x3),
    .io_s(m_1025_io_s),
    .io_cout(m_1025_io_cout)
  );
  Adder m_1026 ( // @[MUL.scala 102:19]
    .io_x1(m_1026_io_x1),
    .io_x2(m_1026_io_x2),
    .io_x3(m_1026_io_x3),
    .io_s(m_1026_io_s),
    .io_cout(m_1026_io_cout)
  );
  Adder m_1027 ( // @[MUL.scala 102:19]
    .io_x1(m_1027_io_x1),
    .io_x2(m_1027_io_x2),
    .io_x3(m_1027_io_x3),
    .io_s(m_1027_io_s),
    .io_cout(m_1027_io_cout)
  );
  Adder m_1028 ( // @[MUL.scala 102:19]
    .io_x1(m_1028_io_x1),
    .io_x2(m_1028_io_x2),
    .io_x3(m_1028_io_x3),
    .io_s(m_1028_io_s),
    .io_cout(m_1028_io_cout)
  );
  Adder m_1029 ( // @[MUL.scala 102:19]
    .io_x1(m_1029_io_x1),
    .io_x2(m_1029_io_x2),
    .io_x3(m_1029_io_x3),
    .io_s(m_1029_io_s),
    .io_cout(m_1029_io_cout)
  );
  Adder m_1030 ( // @[MUL.scala 102:19]
    .io_x1(m_1030_io_x1),
    .io_x2(m_1030_io_x2),
    .io_x3(m_1030_io_x3),
    .io_s(m_1030_io_s),
    .io_cout(m_1030_io_cout)
  );
  Adder m_1031 ( // @[MUL.scala 102:19]
    .io_x1(m_1031_io_x1),
    .io_x2(m_1031_io_x2),
    .io_x3(m_1031_io_x3),
    .io_s(m_1031_io_s),
    .io_cout(m_1031_io_cout)
  );
  Adder m_1032 ( // @[MUL.scala 102:19]
    .io_x1(m_1032_io_x1),
    .io_x2(m_1032_io_x2),
    .io_x3(m_1032_io_x3),
    .io_s(m_1032_io_s),
    .io_cout(m_1032_io_cout)
  );
  Adder m_1033 ( // @[MUL.scala 102:19]
    .io_x1(m_1033_io_x1),
    .io_x2(m_1033_io_x2),
    .io_x3(m_1033_io_x3),
    .io_s(m_1033_io_s),
    .io_cout(m_1033_io_cout)
  );
  Adder m_1034 ( // @[MUL.scala 102:19]
    .io_x1(m_1034_io_x1),
    .io_x2(m_1034_io_x2),
    .io_x3(m_1034_io_x3),
    .io_s(m_1034_io_s),
    .io_cout(m_1034_io_cout)
  );
  Adder m_1035 ( // @[MUL.scala 102:19]
    .io_x1(m_1035_io_x1),
    .io_x2(m_1035_io_x2),
    .io_x3(m_1035_io_x3),
    .io_s(m_1035_io_s),
    .io_cout(m_1035_io_cout)
  );
  Adder m_1036 ( // @[MUL.scala 102:19]
    .io_x1(m_1036_io_x1),
    .io_x2(m_1036_io_x2),
    .io_x3(m_1036_io_x3),
    .io_s(m_1036_io_s),
    .io_cout(m_1036_io_cout)
  );
  Adder m_1037 ( // @[MUL.scala 102:19]
    .io_x1(m_1037_io_x1),
    .io_x2(m_1037_io_x2),
    .io_x3(m_1037_io_x3),
    .io_s(m_1037_io_s),
    .io_cout(m_1037_io_cout)
  );
  Adder m_1038 ( // @[MUL.scala 102:19]
    .io_x1(m_1038_io_x1),
    .io_x2(m_1038_io_x2),
    .io_x3(m_1038_io_x3),
    .io_s(m_1038_io_s),
    .io_cout(m_1038_io_cout)
  );
  Adder m_1039 ( // @[MUL.scala 102:19]
    .io_x1(m_1039_io_x1),
    .io_x2(m_1039_io_x2),
    .io_x3(m_1039_io_x3),
    .io_s(m_1039_io_s),
    .io_cout(m_1039_io_cout)
  );
  Adder m_1040 ( // @[MUL.scala 102:19]
    .io_x1(m_1040_io_x1),
    .io_x2(m_1040_io_x2),
    .io_x3(m_1040_io_x3),
    .io_s(m_1040_io_s),
    .io_cout(m_1040_io_cout)
  );
  Adder m_1041 ( // @[MUL.scala 102:19]
    .io_x1(m_1041_io_x1),
    .io_x2(m_1041_io_x2),
    .io_x3(m_1041_io_x3),
    .io_s(m_1041_io_s),
    .io_cout(m_1041_io_cout)
  );
  Adder m_1042 ( // @[MUL.scala 102:19]
    .io_x1(m_1042_io_x1),
    .io_x2(m_1042_io_x2),
    .io_x3(m_1042_io_x3),
    .io_s(m_1042_io_s),
    .io_cout(m_1042_io_cout)
  );
  Adder m_1043 ( // @[MUL.scala 102:19]
    .io_x1(m_1043_io_x1),
    .io_x2(m_1043_io_x2),
    .io_x3(m_1043_io_x3),
    .io_s(m_1043_io_s),
    .io_cout(m_1043_io_cout)
  );
  Adder m_1044 ( // @[MUL.scala 102:19]
    .io_x1(m_1044_io_x1),
    .io_x2(m_1044_io_x2),
    .io_x3(m_1044_io_x3),
    .io_s(m_1044_io_s),
    .io_cout(m_1044_io_cout)
  );
  Adder m_1045 ( // @[MUL.scala 102:19]
    .io_x1(m_1045_io_x1),
    .io_x2(m_1045_io_x2),
    .io_x3(m_1045_io_x3),
    .io_s(m_1045_io_s),
    .io_cout(m_1045_io_cout)
  );
  Adder m_1046 ( // @[MUL.scala 102:19]
    .io_x1(m_1046_io_x1),
    .io_x2(m_1046_io_x2),
    .io_x3(m_1046_io_x3),
    .io_s(m_1046_io_s),
    .io_cout(m_1046_io_cout)
  );
  Adder m_1047 ( // @[MUL.scala 102:19]
    .io_x1(m_1047_io_x1),
    .io_x2(m_1047_io_x2),
    .io_x3(m_1047_io_x3),
    .io_s(m_1047_io_s),
    .io_cout(m_1047_io_cout)
  );
  Adder m_1048 ( // @[MUL.scala 102:19]
    .io_x1(m_1048_io_x1),
    .io_x2(m_1048_io_x2),
    .io_x3(m_1048_io_x3),
    .io_s(m_1048_io_s),
    .io_cout(m_1048_io_cout)
  );
  Adder m_1049 ( // @[MUL.scala 102:19]
    .io_x1(m_1049_io_x1),
    .io_x2(m_1049_io_x2),
    .io_x3(m_1049_io_x3),
    .io_s(m_1049_io_s),
    .io_cout(m_1049_io_cout)
  );
  Adder m_1050 ( // @[MUL.scala 102:19]
    .io_x1(m_1050_io_x1),
    .io_x2(m_1050_io_x2),
    .io_x3(m_1050_io_x3),
    .io_s(m_1050_io_s),
    .io_cout(m_1050_io_cout)
  );
  Adder m_1051 ( // @[MUL.scala 102:19]
    .io_x1(m_1051_io_x1),
    .io_x2(m_1051_io_x2),
    .io_x3(m_1051_io_x3),
    .io_s(m_1051_io_s),
    .io_cout(m_1051_io_cout)
  );
  Adder m_1052 ( // @[MUL.scala 102:19]
    .io_x1(m_1052_io_x1),
    .io_x2(m_1052_io_x2),
    .io_x3(m_1052_io_x3),
    .io_s(m_1052_io_s),
    .io_cout(m_1052_io_cout)
  );
  Adder m_1053 ( // @[MUL.scala 102:19]
    .io_x1(m_1053_io_x1),
    .io_x2(m_1053_io_x2),
    .io_x3(m_1053_io_x3),
    .io_s(m_1053_io_s),
    .io_cout(m_1053_io_cout)
  );
  Adder m_1054 ( // @[MUL.scala 102:19]
    .io_x1(m_1054_io_x1),
    .io_x2(m_1054_io_x2),
    .io_x3(m_1054_io_x3),
    .io_s(m_1054_io_s),
    .io_cout(m_1054_io_cout)
  );
  Adder m_1055 ( // @[MUL.scala 102:19]
    .io_x1(m_1055_io_x1),
    .io_x2(m_1055_io_x2),
    .io_x3(m_1055_io_x3),
    .io_s(m_1055_io_s),
    .io_cout(m_1055_io_cout)
  );
  Adder m_1056 ( // @[MUL.scala 102:19]
    .io_x1(m_1056_io_x1),
    .io_x2(m_1056_io_x2),
    .io_x3(m_1056_io_x3),
    .io_s(m_1056_io_s),
    .io_cout(m_1056_io_cout)
  );
  Adder m_1057 ( // @[MUL.scala 102:19]
    .io_x1(m_1057_io_x1),
    .io_x2(m_1057_io_x2),
    .io_x3(m_1057_io_x3),
    .io_s(m_1057_io_s),
    .io_cout(m_1057_io_cout)
  );
  Adder m_1058 ( // @[MUL.scala 102:19]
    .io_x1(m_1058_io_x1),
    .io_x2(m_1058_io_x2),
    .io_x3(m_1058_io_x3),
    .io_s(m_1058_io_s),
    .io_cout(m_1058_io_cout)
  );
  Adder m_1059 ( // @[MUL.scala 102:19]
    .io_x1(m_1059_io_x1),
    .io_x2(m_1059_io_x2),
    .io_x3(m_1059_io_x3),
    .io_s(m_1059_io_s),
    .io_cout(m_1059_io_cout)
  );
  Adder m_1060 ( // @[MUL.scala 102:19]
    .io_x1(m_1060_io_x1),
    .io_x2(m_1060_io_x2),
    .io_x3(m_1060_io_x3),
    .io_s(m_1060_io_s),
    .io_cout(m_1060_io_cout)
  );
  Adder m_1061 ( // @[MUL.scala 102:19]
    .io_x1(m_1061_io_x1),
    .io_x2(m_1061_io_x2),
    .io_x3(m_1061_io_x3),
    .io_s(m_1061_io_s),
    .io_cout(m_1061_io_cout)
  );
  Adder m_1062 ( // @[MUL.scala 102:19]
    .io_x1(m_1062_io_x1),
    .io_x2(m_1062_io_x2),
    .io_x3(m_1062_io_x3),
    .io_s(m_1062_io_s),
    .io_cout(m_1062_io_cout)
  );
  Adder m_1063 ( // @[MUL.scala 102:19]
    .io_x1(m_1063_io_x1),
    .io_x2(m_1063_io_x2),
    .io_x3(m_1063_io_x3),
    .io_s(m_1063_io_s),
    .io_cout(m_1063_io_cout)
  );
  Adder m_1064 ( // @[MUL.scala 102:19]
    .io_x1(m_1064_io_x1),
    .io_x2(m_1064_io_x2),
    .io_x3(m_1064_io_x3),
    .io_s(m_1064_io_s),
    .io_cout(m_1064_io_cout)
  );
  Adder m_1065 ( // @[MUL.scala 102:19]
    .io_x1(m_1065_io_x1),
    .io_x2(m_1065_io_x2),
    .io_x3(m_1065_io_x3),
    .io_s(m_1065_io_s),
    .io_cout(m_1065_io_cout)
  );
  Adder m_1066 ( // @[MUL.scala 102:19]
    .io_x1(m_1066_io_x1),
    .io_x2(m_1066_io_x2),
    .io_x3(m_1066_io_x3),
    .io_s(m_1066_io_s),
    .io_cout(m_1066_io_cout)
  );
  Adder m_1067 ( // @[MUL.scala 102:19]
    .io_x1(m_1067_io_x1),
    .io_x2(m_1067_io_x2),
    .io_x3(m_1067_io_x3),
    .io_s(m_1067_io_s),
    .io_cout(m_1067_io_cout)
  );
  Adder m_1068 ( // @[MUL.scala 102:19]
    .io_x1(m_1068_io_x1),
    .io_x2(m_1068_io_x2),
    .io_x3(m_1068_io_x3),
    .io_s(m_1068_io_s),
    .io_cout(m_1068_io_cout)
  );
  Adder m_1069 ( // @[MUL.scala 102:19]
    .io_x1(m_1069_io_x1),
    .io_x2(m_1069_io_x2),
    .io_x3(m_1069_io_x3),
    .io_s(m_1069_io_s),
    .io_cout(m_1069_io_cout)
  );
  Adder m_1070 ( // @[MUL.scala 102:19]
    .io_x1(m_1070_io_x1),
    .io_x2(m_1070_io_x2),
    .io_x3(m_1070_io_x3),
    .io_s(m_1070_io_s),
    .io_cout(m_1070_io_cout)
  );
  Adder m_1071 ( // @[MUL.scala 102:19]
    .io_x1(m_1071_io_x1),
    .io_x2(m_1071_io_x2),
    .io_x3(m_1071_io_x3),
    .io_s(m_1071_io_s),
    .io_cout(m_1071_io_cout)
  );
  Adder m_1072 ( // @[MUL.scala 102:19]
    .io_x1(m_1072_io_x1),
    .io_x2(m_1072_io_x2),
    .io_x3(m_1072_io_x3),
    .io_s(m_1072_io_s),
    .io_cout(m_1072_io_cout)
  );
  Adder m_1073 ( // @[MUL.scala 102:19]
    .io_x1(m_1073_io_x1),
    .io_x2(m_1073_io_x2),
    .io_x3(m_1073_io_x3),
    .io_s(m_1073_io_s),
    .io_cout(m_1073_io_cout)
  );
  Adder m_1074 ( // @[MUL.scala 102:19]
    .io_x1(m_1074_io_x1),
    .io_x2(m_1074_io_x2),
    .io_x3(m_1074_io_x3),
    .io_s(m_1074_io_s),
    .io_cout(m_1074_io_cout)
  );
  Adder m_1075 ( // @[MUL.scala 102:19]
    .io_x1(m_1075_io_x1),
    .io_x2(m_1075_io_x2),
    .io_x3(m_1075_io_x3),
    .io_s(m_1075_io_s),
    .io_cout(m_1075_io_cout)
  );
  Adder m_1076 ( // @[MUL.scala 102:19]
    .io_x1(m_1076_io_x1),
    .io_x2(m_1076_io_x2),
    .io_x3(m_1076_io_x3),
    .io_s(m_1076_io_s),
    .io_cout(m_1076_io_cout)
  );
  Adder m_1077 ( // @[MUL.scala 102:19]
    .io_x1(m_1077_io_x1),
    .io_x2(m_1077_io_x2),
    .io_x3(m_1077_io_x3),
    .io_s(m_1077_io_s),
    .io_cout(m_1077_io_cout)
  );
  Adder m_1078 ( // @[MUL.scala 102:19]
    .io_x1(m_1078_io_x1),
    .io_x2(m_1078_io_x2),
    .io_x3(m_1078_io_x3),
    .io_s(m_1078_io_s),
    .io_cout(m_1078_io_cout)
  );
  Adder m_1079 ( // @[MUL.scala 102:19]
    .io_x1(m_1079_io_x1),
    .io_x2(m_1079_io_x2),
    .io_x3(m_1079_io_x3),
    .io_s(m_1079_io_s),
    .io_cout(m_1079_io_cout)
  );
  Adder m_1080 ( // @[MUL.scala 102:19]
    .io_x1(m_1080_io_x1),
    .io_x2(m_1080_io_x2),
    .io_x3(m_1080_io_x3),
    .io_s(m_1080_io_s),
    .io_cout(m_1080_io_cout)
  );
  Adder m_1081 ( // @[MUL.scala 102:19]
    .io_x1(m_1081_io_x1),
    .io_x2(m_1081_io_x2),
    .io_x3(m_1081_io_x3),
    .io_s(m_1081_io_s),
    .io_cout(m_1081_io_cout)
  );
  Adder m_1082 ( // @[MUL.scala 102:19]
    .io_x1(m_1082_io_x1),
    .io_x2(m_1082_io_x2),
    .io_x3(m_1082_io_x3),
    .io_s(m_1082_io_s),
    .io_cout(m_1082_io_cout)
  );
  Adder m_1083 ( // @[MUL.scala 102:19]
    .io_x1(m_1083_io_x1),
    .io_x2(m_1083_io_x2),
    .io_x3(m_1083_io_x3),
    .io_s(m_1083_io_s),
    .io_cout(m_1083_io_cout)
  );
  Adder m_1084 ( // @[MUL.scala 102:19]
    .io_x1(m_1084_io_x1),
    .io_x2(m_1084_io_x2),
    .io_x3(m_1084_io_x3),
    .io_s(m_1084_io_s),
    .io_cout(m_1084_io_cout)
  );
  Adder m_1085 ( // @[MUL.scala 102:19]
    .io_x1(m_1085_io_x1),
    .io_x2(m_1085_io_x2),
    .io_x3(m_1085_io_x3),
    .io_s(m_1085_io_s),
    .io_cout(m_1085_io_cout)
  );
  Adder m_1086 ( // @[MUL.scala 102:19]
    .io_x1(m_1086_io_x1),
    .io_x2(m_1086_io_x2),
    .io_x3(m_1086_io_x3),
    .io_s(m_1086_io_s),
    .io_cout(m_1086_io_cout)
  );
  Adder m_1087 ( // @[MUL.scala 102:19]
    .io_x1(m_1087_io_x1),
    .io_x2(m_1087_io_x2),
    .io_x3(m_1087_io_x3),
    .io_s(m_1087_io_s),
    .io_cout(m_1087_io_cout)
  );
  Adder m_1088 ( // @[MUL.scala 102:19]
    .io_x1(m_1088_io_x1),
    .io_x2(m_1088_io_x2),
    .io_x3(m_1088_io_x3),
    .io_s(m_1088_io_s),
    .io_cout(m_1088_io_cout)
  );
  Adder m_1089 ( // @[MUL.scala 102:19]
    .io_x1(m_1089_io_x1),
    .io_x2(m_1089_io_x2),
    .io_x3(m_1089_io_x3),
    .io_s(m_1089_io_s),
    .io_cout(m_1089_io_cout)
  );
  Adder m_1090 ( // @[MUL.scala 102:19]
    .io_x1(m_1090_io_x1),
    .io_x2(m_1090_io_x2),
    .io_x3(m_1090_io_x3),
    .io_s(m_1090_io_s),
    .io_cout(m_1090_io_cout)
  );
  Adder m_1091 ( // @[MUL.scala 102:19]
    .io_x1(m_1091_io_x1),
    .io_x2(m_1091_io_x2),
    .io_x3(m_1091_io_x3),
    .io_s(m_1091_io_s),
    .io_cout(m_1091_io_cout)
  );
  Adder m_1092 ( // @[MUL.scala 102:19]
    .io_x1(m_1092_io_x1),
    .io_x2(m_1092_io_x2),
    .io_x3(m_1092_io_x3),
    .io_s(m_1092_io_s),
    .io_cout(m_1092_io_cout)
  );
  Adder m_1093 ( // @[MUL.scala 102:19]
    .io_x1(m_1093_io_x1),
    .io_x2(m_1093_io_x2),
    .io_x3(m_1093_io_x3),
    .io_s(m_1093_io_s),
    .io_cout(m_1093_io_cout)
  );
  Adder m_1094 ( // @[MUL.scala 102:19]
    .io_x1(m_1094_io_x1),
    .io_x2(m_1094_io_x2),
    .io_x3(m_1094_io_x3),
    .io_s(m_1094_io_s),
    .io_cout(m_1094_io_cout)
  );
  Adder m_1095 ( // @[MUL.scala 102:19]
    .io_x1(m_1095_io_x1),
    .io_x2(m_1095_io_x2),
    .io_x3(m_1095_io_x3),
    .io_s(m_1095_io_s),
    .io_cout(m_1095_io_cout)
  );
  Adder m_1096 ( // @[MUL.scala 102:19]
    .io_x1(m_1096_io_x1),
    .io_x2(m_1096_io_x2),
    .io_x3(m_1096_io_x3),
    .io_s(m_1096_io_s),
    .io_cout(m_1096_io_cout)
  );
  Adder m_1097 ( // @[MUL.scala 102:19]
    .io_x1(m_1097_io_x1),
    .io_x2(m_1097_io_x2),
    .io_x3(m_1097_io_x3),
    .io_s(m_1097_io_s),
    .io_cout(m_1097_io_cout)
  );
  Adder m_1098 ( // @[MUL.scala 102:19]
    .io_x1(m_1098_io_x1),
    .io_x2(m_1098_io_x2),
    .io_x3(m_1098_io_x3),
    .io_s(m_1098_io_s),
    .io_cout(m_1098_io_cout)
  );
  Adder m_1099 ( // @[MUL.scala 102:19]
    .io_x1(m_1099_io_x1),
    .io_x2(m_1099_io_x2),
    .io_x3(m_1099_io_x3),
    .io_s(m_1099_io_s),
    .io_cout(m_1099_io_cout)
  );
  Adder m_1100 ( // @[MUL.scala 102:19]
    .io_x1(m_1100_io_x1),
    .io_x2(m_1100_io_x2),
    .io_x3(m_1100_io_x3),
    .io_s(m_1100_io_s),
    .io_cout(m_1100_io_cout)
  );
  Adder m_1101 ( // @[MUL.scala 102:19]
    .io_x1(m_1101_io_x1),
    .io_x2(m_1101_io_x2),
    .io_x3(m_1101_io_x3),
    .io_s(m_1101_io_s),
    .io_cout(m_1101_io_cout)
  );
  Adder m_1102 ( // @[MUL.scala 102:19]
    .io_x1(m_1102_io_x1),
    .io_x2(m_1102_io_x2),
    .io_x3(m_1102_io_x3),
    .io_s(m_1102_io_s),
    .io_cout(m_1102_io_cout)
  );
  Adder m_1103 ( // @[MUL.scala 102:19]
    .io_x1(m_1103_io_x1),
    .io_x2(m_1103_io_x2),
    .io_x3(m_1103_io_x3),
    .io_s(m_1103_io_s),
    .io_cout(m_1103_io_cout)
  );
  Adder m_1104 ( // @[MUL.scala 102:19]
    .io_x1(m_1104_io_x1),
    .io_x2(m_1104_io_x2),
    .io_x3(m_1104_io_x3),
    .io_s(m_1104_io_s),
    .io_cout(m_1104_io_cout)
  );
  Adder m_1105 ( // @[MUL.scala 102:19]
    .io_x1(m_1105_io_x1),
    .io_x2(m_1105_io_x2),
    .io_x3(m_1105_io_x3),
    .io_s(m_1105_io_s),
    .io_cout(m_1105_io_cout)
  );
  Adder m_1106 ( // @[MUL.scala 102:19]
    .io_x1(m_1106_io_x1),
    .io_x2(m_1106_io_x2),
    .io_x3(m_1106_io_x3),
    .io_s(m_1106_io_s),
    .io_cout(m_1106_io_cout)
  );
  Adder m_1107 ( // @[MUL.scala 102:19]
    .io_x1(m_1107_io_x1),
    .io_x2(m_1107_io_x2),
    .io_x3(m_1107_io_x3),
    .io_s(m_1107_io_s),
    .io_cout(m_1107_io_cout)
  );
  Adder m_1108 ( // @[MUL.scala 102:19]
    .io_x1(m_1108_io_x1),
    .io_x2(m_1108_io_x2),
    .io_x3(m_1108_io_x3),
    .io_s(m_1108_io_s),
    .io_cout(m_1108_io_cout)
  );
  Adder m_1109 ( // @[MUL.scala 102:19]
    .io_x1(m_1109_io_x1),
    .io_x2(m_1109_io_x2),
    .io_x3(m_1109_io_x3),
    .io_s(m_1109_io_s),
    .io_cout(m_1109_io_cout)
  );
  Adder m_1110 ( // @[MUL.scala 102:19]
    .io_x1(m_1110_io_x1),
    .io_x2(m_1110_io_x2),
    .io_x3(m_1110_io_x3),
    .io_s(m_1110_io_s),
    .io_cout(m_1110_io_cout)
  );
  Adder m_1111 ( // @[MUL.scala 102:19]
    .io_x1(m_1111_io_x1),
    .io_x2(m_1111_io_x2),
    .io_x3(m_1111_io_x3),
    .io_s(m_1111_io_s),
    .io_cout(m_1111_io_cout)
  );
  Adder m_1112 ( // @[MUL.scala 102:19]
    .io_x1(m_1112_io_x1),
    .io_x2(m_1112_io_x2),
    .io_x3(m_1112_io_x3),
    .io_s(m_1112_io_s),
    .io_cout(m_1112_io_cout)
  );
  Adder m_1113 ( // @[MUL.scala 102:19]
    .io_x1(m_1113_io_x1),
    .io_x2(m_1113_io_x2),
    .io_x3(m_1113_io_x3),
    .io_s(m_1113_io_s),
    .io_cout(m_1113_io_cout)
  );
  Adder m_1114 ( // @[MUL.scala 102:19]
    .io_x1(m_1114_io_x1),
    .io_x2(m_1114_io_x2),
    .io_x3(m_1114_io_x3),
    .io_s(m_1114_io_s),
    .io_cout(m_1114_io_cout)
  );
  Adder m_1115 ( // @[MUL.scala 102:19]
    .io_x1(m_1115_io_x1),
    .io_x2(m_1115_io_x2),
    .io_x3(m_1115_io_x3),
    .io_s(m_1115_io_s),
    .io_cout(m_1115_io_cout)
  );
  Adder m_1116 ( // @[MUL.scala 102:19]
    .io_x1(m_1116_io_x1),
    .io_x2(m_1116_io_x2),
    .io_x3(m_1116_io_x3),
    .io_s(m_1116_io_s),
    .io_cout(m_1116_io_cout)
  );
  Half_Adder m_1117 ( // @[MUL.scala 124:19]
    .io_in_0(m_1117_io_in_0),
    .io_in_1(m_1117_io_in_1),
    .io_out_0(m_1117_io_out_0),
    .io_out_1(m_1117_io_out_1)
  );
  Adder m_1118 ( // @[MUL.scala 102:19]
    .io_x1(m_1118_io_x1),
    .io_x2(m_1118_io_x2),
    .io_x3(m_1118_io_x3),
    .io_s(m_1118_io_s),
    .io_cout(m_1118_io_cout)
  );
  Adder m_1119 ( // @[MUL.scala 102:19]
    .io_x1(m_1119_io_x1),
    .io_x2(m_1119_io_x2),
    .io_x3(m_1119_io_x3),
    .io_s(m_1119_io_s),
    .io_cout(m_1119_io_cout)
  );
  Adder m_1120 ( // @[MUL.scala 102:19]
    .io_x1(m_1120_io_x1),
    .io_x2(m_1120_io_x2),
    .io_x3(m_1120_io_x3),
    .io_s(m_1120_io_s),
    .io_cout(m_1120_io_cout)
  );
  Adder m_1121 ( // @[MUL.scala 102:19]
    .io_x1(m_1121_io_x1),
    .io_x2(m_1121_io_x2),
    .io_x3(m_1121_io_x3),
    .io_s(m_1121_io_s),
    .io_cout(m_1121_io_cout)
  );
  Adder m_1122 ( // @[MUL.scala 102:19]
    .io_x1(m_1122_io_x1),
    .io_x2(m_1122_io_x2),
    .io_x3(m_1122_io_x3),
    .io_s(m_1122_io_s),
    .io_cout(m_1122_io_cout)
  );
  Adder m_1123 ( // @[MUL.scala 102:19]
    .io_x1(m_1123_io_x1),
    .io_x2(m_1123_io_x2),
    .io_x3(m_1123_io_x3),
    .io_s(m_1123_io_s),
    .io_cout(m_1123_io_cout)
  );
  Half_Adder m_1124 ( // @[MUL.scala 124:19]
    .io_in_0(m_1124_io_in_0),
    .io_in_1(m_1124_io_in_1),
    .io_out_0(m_1124_io_out_0),
    .io_out_1(m_1124_io_out_1)
  );
  Adder m_1125 ( // @[MUL.scala 102:19]
    .io_x1(m_1125_io_x1),
    .io_x2(m_1125_io_x2),
    .io_x3(m_1125_io_x3),
    .io_s(m_1125_io_s),
    .io_cout(m_1125_io_cout)
  );
  Adder m_1126 ( // @[MUL.scala 102:19]
    .io_x1(m_1126_io_x1),
    .io_x2(m_1126_io_x2),
    .io_x3(m_1126_io_x3),
    .io_s(m_1126_io_s),
    .io_cout(m_1126_io_cout)
  );
  Adder m_1127 ( // @[MUL.scala 102:19]
    .io_x1(m_1127_io_x1),
    .io_x2(m_1127_io_x2),
    .io_x3(m_1127_io_x3),
    .io_s(m_1127_io_s),
    .io_cout(m_1127_io_cout)
  );
  Adder m_1128 ( // @[MUL.scala 102:19]
    .io_x1(m_1128_io_x1),
    .io_x2(m_1128_io_x2),
    .io_x3(m_1128_io_x3),
    .io_s(m_1128_io_s),
    .io_cout(m_1128_io_cout)
  );
  Adder m_1129 ( // @[MUL.scala 102:19]
    .io_x1(m_1129_io_x1),
    .io_x2(m_1129_io_x2),
    .io_x3(m_1129_io_x3),
    .io_s(m_1129_io_s),
    .io_cout(m_1129_io_cout)
  );
  Adder m_1130 ( // @[MUL.scala 102:19]
    .io_x1(m_1130_io_x1),
    .io_x2(m_1130_io_x2),
    .io_x3(m_1130_io_x3),
    .io_s(m_1130_io_s),
    .io_cout(m_1130_io_cout)
  );
  Half_Adder m_1131 ( // @[MUL.scala 124:19]
    .io_in_0(m_1131_io_in_0),
    .io_in_1(m_1131_io_in_1),
    .io_out_0(m_1131_io_out_0),
    .io_out_1(m_1131_io_out_1)
  );
  Adder m_1132 ( // @[MUL.scala 102:19]
    .io_x1(m_1132_io_x1),
    .io_x2(m_1132_io_x2),
    .io_x3(m_1132_io_x3),
    .io_s(m_1132_io_s),
    .io_cout(m_1132_io_cout)
  );
  Adder m_1133 ( // @[MUL.scala 102:19]
    .io_x1(m_1133_io_x1),
    .io_x2(m_1133_io_x2),
    .io_x3(m_1133_io_x3),
    .io_s(m_1133_io_s),
    .io_cout(m_1133_io_cout)
  );
  Adder m_1134 ( // @[MUL.scala 102:19]
    .io_x1(m_1134_io_x1),
    .io_x2(m_1134_io_x2),
    .io_x3(m_1134_io_x3),
    .io_s(m_1134_io_s),
    .io_cout(m_1134_io_cout)
  );
  Adder m_1135 ( // @[MUL.scala 102:19]
    .io_x1(m_1135_io_x1),
    .io_x2(m_1135_io_x2),
    .io_x3(m_1135_io_x3),
    .io_s(m_1135_io_s),
    .io_cout(m_1135_io_cout)
  );
  Adder m_1136 ( // @[MUL.scala 102:19]
    .io_x1(m_1136_io_x1),
    .io_x2(m_1136_io_x2),
    .io_x3(m_1136_io_x3),
    .io_s(m_1136_io_s),
    .io_cout(m_1136_io_cout)
  );
  Adder m_1137 ( // @[MUL.scala 102:19]
    .io_x1(m_1137_io_x1),
    .io_x2(m_1137_io_x2),
    .io_x3(m_1137_io_x3),
    .io_s(m_1137_io_s),
    .io_cout(m_1137_io_cout)
  );
  Half_Adder m_1138 ( // @[MUL.scala 124:19]
    .io_in_0(m_1138_io_in_0),
    .io_in_1(m_1138_io_in_1),
    .io_out_0(m_1138_io_out_0),
    .io_out_1(m_1138_io_out_1)
  );
  Adder m_1139 ( // @[MUL.scala 102:19]
    .io_x1(m_1139_io_x1),
    .io_x2(m_1139_io_x2),
    .io_x3(m_1139_io_x3),
    .io_s(m_1139_io_s),
    .io_cout(m_1139_io_cout)
  );
  Adder m_1140 ( // @[MUL.scala 102:19]
    .io_x1(m_1140_io_x1),
    .io_x2(m_1140_io_x2),
    .io_x3(m_1140_io_x3),
    .io_s(m_1140_io_s),
    .io_cout(m_1140_io_cout)
  );
  Adder m_1141 ( // @[MUL.scala 102:19]
    .io_x1(m_1141_io_x1),
    .io_x2(m_1141_io_x2),
    .io_x3(m_1141_io_x3),
    .io_s(m_1141_io_s),
    .io_cout(m_1141_io_cout)
  );
  Adder m_1142 ( // @[MUL.scala 102:19]
    .io_x1(m_1142_io_x1),
    .io_x2(m_1142_io_x2),
    .io_x3(m_1142_io_x3),
    .io_s(m_1142_io_s),
    .io_cout(m_1142_io_cout)
  );
  Adder m_1143 ( // @[MUL.scala 102:19]
    .io_x1(m_1143_io_x1),
    .io_x2(m_1143_io_x2),
    .io_x3(m_1143_io_x3),
    .io_s(m_1143_io_s),
    .io_cout(m_1143_io_cout)
  );
  Adder m_1144 ( // @[MUL.scala 102:19]
    .io_x1(m_1144_io_x1),
    .io_x2(m_1144_io_x2),
    .io_x3(m_1144_io_x3),
    .io_s(m_1144_io_s),
    .io_cout(m_1144_io_cout)
  );
  Half_Adder m_1145 ( // @[MUL.scala 124:19]
    .io_in_0(m_1145_io_in_0),
    .io_in_1(m_1145_io_in_1),
    .io_out_0(m_1145_io_out_0),
    .io_out_1(m_1145_io_out_1)
  );
  Adder m_1146 ( // @[MUL.scala 102:19]
    .io_x1(m_1146_io_x1),
    .io_x2(m_1146_io_x2),
    .io_x3(m_1146_io_x3),
    .io_s(m_1146_io_s),
    .io_cout(m_1146_io_cout)
  );
  Adder m_1147 ( // @[MUL.scala 102:19]
    .io_x1(m_1147_io_x1),
    .io_x2(m_1147_io_x2),
    .io_x3(m_1147_io_x3),
    .io_s(m_1147_io_s),
    .io_cout(m_1147_io_cout)
  );
  Adder m_1148 ( // @[MUL.scala 102:19]
    .io_x1(m_1148_io_x1),
    .io_x2(m_1148_io_x2),
    .io_x3(m_1148_io_x3),
    .io_s(m_1148_io_s),
    .io_cout(m_1148_io_cout)
  );
  Adder m_1149 ( // @[MUL.scala 102:19]
    .io_x1(m_1149_io_x1),
    .io_x2(m_1149_io_x2),
    .io_x3(m_1149_io_x3),
    .io_s(m_1149_io_s),
    .io_cout(m_1149_io_cout)
  );
  Adder m_1150 ( // @[MUL.scala 102:19]
    .io_x1(m_1150_io_x1),
    .io_x2(m_1150_io_x2),
    .io_x3(m_1150_io_x3),
    .io_s(m_1150_io_s),
    .io_cout(m_1150_io_cout)
  );
  Adder m_1151 ( // @[MUL.scala 102:19]
    .io_x1(m_1151_io_x1),
    .io_x2(m_1151_io_x2),
    .io_x3(m_1151_io_x3),
    .io_s(m_1151_io_s),
    .io_cout(m_1151_io_cout)
  );
  Adder m_1152 ( // @[MUL.scala 102:19]
    .io_x1(m_1152_io_x1),
    .io_x2(m_1152_io_x2),
    .io_x3(m_1152_io_x3),
    .io_s(m_1152_io_s),
    .io_cout(m_1152_io_cout)
  );
  Adder m_1153 ( // @[MUL.scala 102:19]
    .io_x1(m_1153_io_x1),
    .io_x2(m_1153_io_x2),
    .io_x3(m_1153_io_x3),
    .io_s(m_1153_io_s),
    .io_cout(m_1153_io_cout)
  );
  Adder m_1154 ( // @[MUL.scala 102:19]
    .io_x1(m_1154_io_x1),
    .io_x2(m_1154_io_x2),
    .io_x3(m_1154_io_x3),
    .io_s(m_1154_io_s),
    .io_cout(m_1154_io_cout)
  );
  Adder m_1155 ( // @[MUL.scala 102:19]
    .io_x1(m_1155_io_x1),
    .io_x2(m_1155_io_x2),
    .io_x3(m_1155_io_x3),
    .io_s(m_1155_io_s),
    .io_cout(m_1155_io_cout)
  );
  Adder m_1156 ( // @[MUL.scala 102:19]
    .io_x1(m_1156_io_x1),
    .io_x2(m_1156_io_x2),
    .io_x3(m_1156_io_x3),
    .io_s(m_1156_io_s),
    .io_cout(m_1156_io_cout)
  );
  Adder m_1157 ( // @[MUL.scala 102:19]
    .io_x1(m_1157_io_x1),
    .io_x2(m_1157_io_x2),
    .io_x3(m_1157_io_x3),
    .io_s(m_1157_io_s),
    .io_cout(m_1157_io_cout)
  );
  Adder m_1158 ( // @[MUL.scala 102:19]
    .io_x1(m_1158_io_x1),
    .io_x2(m_1158_io_x2),
    .io_x3(m_1158_io_x3),
    .io_s(m_1158_io_s),
    .io_cout(m_1158_io_cout)
  );
  Adder m_1159 ( // @[MUL.scala 102:19]
    .io_x1(m_1159_io_x1),
    .io_x2(m_1159_io_x2),
    .io_x3(m_1159_io_x3),
    .io_s(m_1159_io_s),
    .io_cout(m_1159_io_cout)
  );
  Adder m_1160 ( // @[MUL.scala 102:19]
    .io_x1(m_1160_io_x1),
    .io_x2(m_1160_io_x2),
    .io_x3(m_1160_io_x3),
    .io_s(m_1160_io_s),
    .io_cout(m_1160_io_cout)
  );
  Adder m_1161 ( // @[MUL.scala 102:19]
    .io_x1(m_1161_io_x1),
    .io_x2(m_1161_io_x2),
    .io_x3(m_1161_io_x3),
    .io_s(m_1161_io_s),
    .io_cout(m_1161_io_cout)
  );
  Adder m_1162 ( // @[MUL.scala 102:19]
    .io_x1(m_1162_io_x1),
    .io_x2(m_1162_io_x2),
    .io_x3(m_1162_io_x3),
    .io_s(m_1162_io_s),
    .io_cout(m_1162_io_cout)
  );
  Adder m_1163 ( // @[MUL.scala 102:19]
    .io_x1(m_1163_io_x1),
    .io_x2(m_1163_io_x2),
    .io_x3(m_1163_io_x3),
    .io_s(m_1163_io_s),
    .io_cout(m_1163_io_cout)
  );
  Adder m_1164 ( // @[MUL.scala 102:19]
    .io_x1(m_1164_io_x1),
    .io_x2(m_1164_io_x2),
    .io_x3(m_1164_io_x3),
    .io_s(m_1164_io_s),
    .io_cout(m_1164_io_cout)
  );
  Adder m_1165 ( // @[MUL.scala 102:19]
    .io_x1(m_1165_io_x1),
    .io_x2(m_1165_io_x2),
    .io_x3(m_1165_io_x3),
    .io_s(m_1165_io_s),
    .io_cout(m_1165_io_cout)
  );
  Adder m_1166 ( // @[MUL.scala 102:19]
    .io_x1(m_1166_io_x1),
    .io_x2(m_1166_io_x2),
    .io_x3(m_1166_io_x3),
    .io_s(m_1166_io_s),
    .io_cout(m_1166_io_cout)
  );
  Adder m_1167 ( // @[MUL.scala 102:19]
    .io_x1(m_1167_io_x1),
    .io_x2(m_1167_io_x2),
    .io_x3(m_1167_io_x3),
    .io_s(m_1167_io_s),
    .io_cout(m_1167_io_cout)
  );
  Adder m_1168 ( // @[MUL.scala 102:19]
    .io_x1(m_1168_io_x1),
    .io_x2(m_1168_io_x2),
    .io_x3(m_1168_io_x3),
    .io_s(m_1168_io_s),
    .io_cout(m_1168_io_cout)
  );
  Adder m_1169 ( // @[MUL.scala 102:19]
    .io_x1(m_1169_io_x1),
    .io_x2(m_1169_io_x2),
    .io_x3(m_1169_io_x3),
    .io_s(m_1169_io_s),
    .io_cout(m_1169_io_cout)
  );
  Adder m_1170 ( // @[MUL.scala 102:19]
    .io_x1(m_1170_io_x1),
    .io_x2(m_1170_io_x2),
    .io_x3(m_1170_io_x3),
    .io_s(m_1170_io_s),
    .io_cout(m_1170_io_cout)
  );
  Adder m_1171 ( // @[MUL.scala 102:19]
    .io_x1(m_1171_io_x1),
    .io_x2(m_1171_io_x2),
    .io_x3(m_1171_io_x3),
    .io_s(m_1171_io_s),
    .io_cout(m_1171_io_cout)
  );
  Adder m_1172 ( // @[MUL.scala 102:19]
    .io_x1(m_1172_io_x1),
    .io_x2(m_1172_io_x2),
    .io_x3(m_1172_io_x3),
    .io_s(m_1172_io_s),
    .io_cout(m_1172_io_cout)
  );
  Adder m_1173 ( // @[MUL.scala 102:19]
    .io_x1(m_1173_io_x1),
    .io_x2(m_1173_io_x2),
    .io_x3(m_1173_io_x3),
    .io_s(m_1173_io_s),
    .io_cout(m_1173_io_cout)
  );
  Adder m_1174 ( // @[MUL.scala 102:19]
    .io_x1(m_1174_io_x1),
    .io_x2(m_1174_io_x2),
    .io_x3(m_1174_io_x3),
    .io_s(m_1174_io_s),
    .io_cout(m_1174_io_cout)
  );
  Adder m_1175 ( // @[MUL.scala 102:19]
    .io_x1(m_1175_io_x1),
    .io_x2(m_1175_io_x2),
    .io_x3(m_1175_io_x3),
    .io_s(m_1175_io_s),
    .io_cout(m_1175_io_cout)
  );
  Adder m_1176 ( // @[MUL.scala 102:19]
    .io_x1(m_1176_io_x1),
    .io_x2(m_1176_io_x2),
    .io_x3(m_1176_io_x3),
    .io_s(m_1176_io_s),
    .io_cout(m_1176_io_cout)
  );
  Adder m_1177 ( // @[MUL.scala 102:19]
    .io_x1(m_1177_io_x1),
    .io_x2(m_1177_io_x2),
    .io_x3(m_1177_io_x3),
    .io_s(m_1177_io_s),
    .io_cout(m_1177_io_cout)
  );
  Adder m_1178 ( // @[MUL.scala 102:19]
    .io_x1(m_1178_io_x1),
    .io_x2(m_1178_io_x2),
    .io_x3(m_1178_io_x3),
    .io_s(m_1178_io_s),
    .io_cout(m_1178_io_cout)
  );
  Adder m_1179 ( // @[MUL.scala 102:19]
    .io_x1(m_1179_io_x1),
    .io_x2(m_1179_io_x2),
    .io_x3(m_1179_io_x3),
    .io_s(m_1179_io_s),
    .io_cout(m_1179_io_cout)
  );
  Adder m_1180 ( // @[MUL.scala 102:19]
    .io_x1(m_1180_io_x1),
    .io_x2(m_1180_io_x2),
    .io_x3(m_1180_io_x3),
    .io_s(m_1180_io_s),
    .io_cout(m_1180_io_cout)
  );
  Adder m_1181 ( // @[MUL.scala 102:19]
    .io_x1(m_1181_io_x1),
    .io_x2(m_1181_io_x2),
    .io_x3(m_1181_io_x3),
    .io_s(m_1181_io_s),
    .io_cout(m_1181_io_cout)
  );
  Adder m_1182 ( // @[MUL.scala 102:19]
    .io_x1(m_1182_io_x1),
    .io_x2(m_1182_io_x2),
    .io_x3(m_1182_io_x3),
    .io_s(m_1182_io_s),
    .io_cout(m_1182_io_cout)
  );
  Adder m_1183 ( // @[MUL.scala 102:19]
    .io_x1(m_1183_io_x1),
    .io_x2(m_1183_io_x2),
    .io_x3(m_1183_io_x3),
    .io_s(m_1183_io_s),
    .io_cout(m_1183_io_cout)
  );
  Adder m_1184 ( // @[MUL.scala 102:19]
    .io_x1(m_1184_io_x1),
    .io_x2(m_1184_io_x2),
    .io_x3(m_1184_io_x3),
    .io_s(m_1184_io_s),
    .io_cout(m_1184_io_cout)
  );
  Adder m_1185 ( // @[MUL.scala 102:19]
    .io_x1(m_1185_io_x1),
    .io_x2(m_1185_io_x2),
    .io_x3(m_1185_io_x3),
    .io_s(m_1185_io_s),
    .io_cout(m_1185_io_cout)
  );
  Adder m_1186 ( // @[MUL.scala 102:19]
    .io_x1(m_1186_io_x1),
    .io_x2(m_1186_io_x2),
    .io_x3(m_1186_io_x3),
    .io_s(m_1186_io_s),
    .io_cout(m_1186_io_cout)
  );
  Half_Adder m_1187 ( // @[MUL.scala 124:19]
    .io_in_0(m_1187_io_in_0),
    .io_in_1(m_1187_io_in_1),
    .io_out_0(m_1187_io_out_0),
    .io_out_1(m_1187_io_out_1)
  );
  Adder m_1188 ( // @[MUL.scala 102:19]
    .io_x1(m_1188_io_x1),
    .io_x2(m_1188_io_x2),
    .io_x3(m_1188_io_x3),
    .io_s(m_1188_io_s),
    .io_cout(m_1188_io_cout)
  );
  Adder m_1189 ( // @[MUL.scala 102:19]
    .io_x1(m_1189_io_x1),
    .io_x2(m_1189_io_x2),
    .io_x3(m_1189_io_x3),
    .io_s(m_1189_io_s),
    .io_cout(m_1189_io_cout)
  );
  Adder m_1190 ( // @[MUL.scala 102:19]
    .io_x1(m_1190_io_x1),
    .io_x2(m_1190_io_x2),
    .io_x3(m_1190_io_x3),
    .io_s(m_1190_io_s),
    .io_cout(m_1190_io_cout)
  );
  Adder m_1191 ( // @[MUL.scala 102:19]
    .io_x1(m_1191_io_x1),
    .io_x2(m_1191_io_x2),
    .io_x3(m_1191_io_x3),
    .io_s(m_1191_io_s),
    .io_cout(m_1191_io_cout)
  );
  Adder m_1192 ( // @[MUL.scala 102:19]
    .io_x1(m_1192_io_x1),
    .io_x2(m_1192_io_x2),
    .io_x3(m_1192_io_x3),
    .io_s(m_1192_io_s),
    .io_cout(m_1192_io_cout)
  );
  Adder m_1193 ( // @[MUL.scala 102:19]
    .io_x1(m_1193_io_x1),
    .io_x2(m_1193_io_x2),
    .io_x3(m_1193_io_x3),
    .io_s(m_1193_io_s),
    .io_cout(m_1193_io_cout)
  );
  Adder m_1194 ( // @[MUL.scala 102:19]
    .io_x1(m_1194_io_x1),
    .io_x2(m_1194_io_x2),
    .io_x3(m_1194_io_x3),
    .io_s(m_1194_io_s),
    .io_cout(m_1194_io_cout)
  );
  Adder m_1195 ( // @[MUL.scala 102:19]
    .io_x1(m_1195_io_x1),
    .io_x2(m_1195_io_x2),
    .io_x3(m_1195_io_x3),
    .io_s(m_1195_io_s),
    .io_cout(m_1195_io_cout)
  );
  Adder m_1196 ( // @[MUL.scala 102:19]
    .io_x1(m_1196_io_x1),
    .io_x2(m_1196_io_x2),
    .io_x3(m_1196_io_x3),
    .io_s(m_1196_io_s),
    .io_cout(m_1196_io_cout)
  );
  Adder m_1197 ( // @[MUL.scala 102:19]
    .io_x1(m_1197_io_x1),
    .io_x2(m_1197_io_x2),
    .io_x3(m_1197_io_x3),
    .io_s(m_1197_io_s),
    .io_cout(m_1197_io_cout)
  );
  Adder m_1198 ( // @[MUL.scala 102:19]
    .io_x1(m_1198_io_x1),
    .io_x2(m_1198_io_x2),
    .io_x3(m_1198_io_x3),
    .io_s(m_1198_io_s),
    .io_cout(m_1198_io_cout)
  );
  Adder m_1199 ( // @[MUL.scala 102:19]
    .io_x1(m_1199_io_x1),
    .io_x2(m_1199_io_x2),
    .io_x3(m_1199_io_x3),
    .io_s(m_1199_io_s),
    .io_cout(m_1199_io_cout)
  );
  Adder m_1200 ( // @[MUL.scala 102:19]
    .io_x1(m_1200_io_x1),
    .io_x2(m_1200_io_x2),
    .io_x3(m_1200_io_x3),
    .io_s(m_1200_io_s),
    .io_cout(m_1200_io_cout)
  );
  Adder m_1201 ( // @[MUL.scala 102:19]
    .io_x1(m_1201_io_x1),
    .io_x2(m_1201_io_x2),
    .io_x3(m_1201_io_x3),
    .io_s(m_1201_io_s),
    .io_cout(m_1201_io_cout)
  );
  Adder m_1202 ( // @[MUL.scala 102:19]
    .io_x1(m_1202_io_x1),
    .io_x2(m_1202_io_x2),
    .io_x3(m_1202_io_x3),
    .io_s(m_1202_io_s),
    .io_cout(m_1202_io_cout)
  );
  Adder m_1203 ( // @[MUL.scala 102:19]
    .io_x1(m_1203_io_x1),
    .io_x2(m_1203_io_x2),
    .io_x3(m_1203_io_x3),
    .io_s(m_1203_io_s),
    .io_cout(m_1203_io_cout)
  );
  Adder m_1204 ( // @[MUL.scala 102:19]
    .io_x1(m_1204_io_x1),
    .io_x2(m_1204_io_x2),
    .io_x3(m_1204_io_x3),
    .io_s(m_1204_io_s),
    .io_cout(m_1204_io_cout)
  );
  Adder m_1205 ( // @[MUL.scala 102:19]
    .io_x1(m_1205_io_x1),
    .io_x2(m_1205_io_x2),
    .io_x3(m_1205_io_x3),
    .io_s(m_1205_io_s),
    .io_cout(m_1205_io_cout)
  );
  Adder m_1206 ( // @[MUL.scala 102:19]
    .io_x1(m_1206_io_x1),
    .io_x2(m_1206_io_x2),
    .io_x3(m_1206_io_x3),
    .io_s(m_1206_io_s),
    .io_cout(m_1206_io_cout)
  );
  Adder m_1207 ( // @[MUL.scala 102:19]
    .io_x1(m_1207_io_x1),
    .io_x2(m_1207_io_x2),
    .io_x3(m_1207_io_x3),
    .io_s(m_1207_io_s),
    .io_cout(m_1207_io_cout)
  );
  Adder m_1208 ( // @[MUL.scala 102:19]
    .io_x1(m_1208_io_x1),
    .io_x2(m_1208_io_x2),
    .io_x3(m_1208_io_x3),
    .io_s(m_1208_io_s),
    .io_cout(m_1208_io_cout)
  );
  Adder m_1209 ( // @[MUL.scala 102:19]
    .io_x1(m_1209_io_x1),
    .io_x2(m_1209_io_x2),
    .io_x3(m_1209_io_x3),
    .io_s(m_1209_io_s),
    .io_cout(m_1209_io_cout)
  );
  Adder m_1210 ( // @[MUL.scala 102:19]
    .io_x1(m_1210_io_x1),
    .io_x2(m_1210_io_x2),
    .io_x3(m_1210_io_x3),
    .io_s(m_1210_io_s),
    .io_cout(m_1210_io_cout)
  );
  Adder m_1211 ( // @[MUL.scala 102:19]
    .io_x1(m_1211_io_x1),
    .io_x2(m_1211_io_x2),
    .io_x3(m_1211_io_x3),
    .io_s(m_1211_io_s),
    .io_cout(m_1211_io_cout)
  );
  Adder m_1212 ( // @[MUL.scala 102:19]
    .io_x1(m_1212_io_x1),
    .io_x2(m_1212_io_x2),
    .io_x3(m_1212_io_x3),
    .io_s(m_1212_io_s),
    .io_cout(m_1212_io_cout)
  );
  Adder m_1213 ( // @[MUL.scala 102:19]
    .io_x1(m_1213_io_x1),
    .io_x2(m_1213_io_x2),
    .io_x3(m_1213_io_x3),
    .io_s(m_1213_io_s),
    .io_cout(m_1213_io_cout)
  );
  Adder m_1214 ( // @[MUL.scala 102:19]
    .io_x1(m_1214_io_x1),
    .io_x2(m_1214_io_x2),
    .io_x3(m_1214_io_x3),
    .io_s(m_1214_io_s),
    .io_cout(m_1214_io_cout)
  );
  Adder m_1215 ( // @[MUL.scala 102:19]
    .io_x1(m_1215_io_x1),
    .io_x2(m_1215_io_x2),
    .io_x3(m_1215_io_x3),
    .io_s(m_1215_io_s),
    .io_cout(m_1215_io_cout)
  );
  Adder m_1216 ( // @[MUL.scala 102:19]
    .io_x1(m_1216_io_x1),
    .io_x2(m_1216_io_x2),
    .io_x3(m_1216_io_x3),
    .io_s(m_1216_io_s),
    .io_cout(m_1216_io_cout)
  );
  Adder m_1217 ( // @[MUL.scala 102:19]
    .io_x1(m_1217_io_x1),
    .io_x2(m_1217_io_x2),
    .io_x3(m_1217_io_x3),
    .io_s(m_1217_io_s),
    .io_cout(m_1217_io_cout)
  );
  Adder m_1218 ( // @[MUL.scala 102:19]
    .io_x1(m_1218_io_x1),
    .io_x2(m_1218_io_x2),
    .io_x3(m_1218_io_x3),
    .io_s(m_1218_io_s),
    .io_cout(m_1218_io_cout)
  );
  Adder m_1219 ( // @[MUL.scala 102:19]
    .io_x1(m_1219_io_x1),
    .io_x2(m_1219_io_x2),
    .io_x3(m_1219_io_x3),
    .io_s(m_1219_io_s),
    .io_cout(m_1219_io_cout)
  );
  Adder m_1220 ( // @[MUL.scala 102:19]
    .io_x1(m_1220_io_x1),
    .io_x2(m_1220_io_x2),
    .io_x3(m_1220_io_x3),
    .io_s(m_1220_io_s),
    .io_cout(m_1220_io_cout)
  );
  Adder m_1221 ( // @[MUL.scala 102:19]
    .io_x1(m_1221_io_x1),
    .io_x2(m_1221_io_x2),
    .io_x3(m_1221_io_x3),
    .io_s(m_1221_io_s),
    .io_cout(m_1221_io_cout)
  );
  Half_Adder m_1222 ( // @[MUL.scala 124:19]
    .io_in_0(m_1222_io_in_0),
    .io_in_1(m_1222_io_in_1),
    .io_out_0(m_1222_io_out_0),
    .io_out_1(m_1222_io_out_1)
  );
  Adder m_1223 ( // @[MUL.scala 102:19]
    .io_x1(m_1223_io_x1),
    .io_x2(m_1223_io_x2),
    .io_x3(m_1223_io_x3),
    .io_s(m_1223_io_s),
    .io_cout(m_1223_io_cout)
  );
  Adder m_1224 ( // @[MUL.scala 102:19]
    .io_x1(m_1224_io_x1),
    .io_x2(m_1224_io_x2),
    .io_x3(m_1224_io_x3),
    .io_s(m_1224_io_s),
    .io_cout(m_1224_io_cout)
  );
  Adder m_1225 ( // @[MUL.scala 102:19]
    .io_x1(m_1225_io_x1),
    .io_x2(m_1225_io_x2),
    .io_x3(m_1225_io_x3),
    .io_s(m_1225_io_s),
    .io_cout(m_1225_io_cout)
  );
  Adder m_1226 ( // @[MUL.scala 102:19]
    .io_x1(m_1226_io_x1),
    .io_x2(m_1226_io_x2),
    .io_x3(m_1226_io_x3),
    .io_s(m_1226_io_s),
    .io_cout(m_1226_io_cout)
  );
  Half_Adder m_1227 ( // @[MUL.scala 124:19]
    .io_in_0(m_1227_io_in_0),
    .io_in_1(m_1227_io_in_1),
    .io_out_0(m_1227_io_out_0),
    .io_out_1(m_1227_io_out_1)
  );
  Adder m_1228 ( // @[MUL.scala 102:19]
    .io_x1(m_1228_io_x1),
    .io_x2(m_1228_io_x2),
    .io_x3(m_1228_io_x3),
    .io_s(m_1228_io_s),
    .io_cout(m_1228_io_cout)
  );
  Adder m_1229 ( // @[MUL.scala 102:19]
    .io_x1(m_1229_io_x1),
    .io_x2(m_1229_io_x2),
    .io_x3(m_1229_io_x3),
    .io_s(m_1229_io_s),
    .io_cout(m_1229_io_cout)
  );
  Adder m_1230 ( // @[MUL.scala 102:19]
    .io_x1(m_1230_io_x1),
    .io_x2(m_1230_io_x2),
    .io_x3(m_1230_io_x3),
    .io_s(m_1230_io_s),
    .io_cout(m_1230_io_cout)
  );
  Adder m_1231 ( // @[MUL.scala 102:19]
    .io_x1(m_1231_io_x1),
    .io_x2(m_1231_io_x2),
    .io_x3(m_1231_io_x3),
    .io_s(m_1231_io_s),
    .io_cout(m_1231_io_cout)
  );
  Half_Adder m_1232 ( // @[MUL.scala 124:19]
    .io_in_0(m_1232_io_in_0),
    .io_in_1(m_1232_io_in_1),
    .io_out_0(m_1232_io_out_0),
    .io_out_1(m_1232_io_out_1)
  );
  Adder m_1233 ( // @[MUL.scala 102:19]
    .io_x1(m_1233_io_x1),
    .io_x2(m_1233_io_x2),
    .io_x3(m_1233_io_x3),
    .io_s(m_1233_io_s),
    .io_cout(m_1233_io_cout)
  );
  Adder m_1234 ( // @[MUL.scala 102:19]
    .io_x1(m_1234_io_x1),
    .io_x2(m_1234_io_x2),
    .io_x3(m_1234_io_x3),
    .io_s(m_1234_io_s),
    .io_cout(m_1234_io_cout)
  );
  Adder m_1235 ( // @[MUL.scala 102:19]
    .io_x1(m_1235_io_x1),
    .io_x2(m_1235_io_x2),
    .io_x3(m_1235_io_x3),
    .io_s(m_1235_io_s),
    .io_cout(m_1235_io_cout)
  );
  Adder m_1236 ( // @[MUL.scala 102:19]
    .io_x1(m_1236_io_x1),
    .io_x2(m_1236_io_x2),
    .io_x3(m_1236_io_x3),
    .io_s(m_1236_io_s),
    .io_cout(m_1236_io_cout)
  );
  Half_Adder m_1237 ( // @[MUL.scala 124:19]
    .io_in_0(m_1237_io_in_0),
    .io_in_1(m_1237_io_in_1),
    .io_out_0(m_1237_io_out_0),
    .io_out_1(m_1237_io_out_1)
  );
  Adder m_1238 ( // @[MUL.scala 102:19]
    .io_x1(m_1238_io_x1),
    .io_x2(m_1238_io_x2),
    .io_x3(m_1238_io_x3),
    .io_s(m_1238_io_s),
    .io_cout(m_1238_io_cout)
  );
  Adder m_1239 ( // @[MUL.scala 102:19]
    .io_x1(m_1239_io_x1),
    .io_x2(m_1239_io_x2),
    .io_x3(m_1239_io_x3),
    .io_s(m_1239_io_s),
    .io_cout(m_1239_io_cout)
  );
  Adder m_1240 ( // @[MUL.scala 102:19]
    .io_x1(m_1240_io_x1),
    .io_x2(m_1240_io_x2),
    .io_x3(m_1240_io_x3),
    .io_s(m_1240_io_s),
    .io_cout(m_1240_io_cout)
  );
  Adder m_1241 ( // @[MUL.scala 102:19]
    .io_x1(m_1241_io_x1),
    .io_x2(m_1241_io_x2),
    .io_x3(m_1241_io_x3),
    .io_s(m_1241_io_s),
    .io_cout(m_1241_io_cout)
  );
  Half_Adder m_1242 ( // @[MUL.scala 124:19]
    .io_in_0(m_1242_io_in_0),
    .io_in_1(m_1242_io_in_1),
    .io_out_0(m_1242_io_out_0),
    .io_out_1(m_1242_io_out_1)
  );
  Adder m_1243 ( // @[MUL.scala 102:19]
    .io_x1(m_1243_io_x1),
    .io_x2(m_1243_io_x2),
    .io_x3(m_1243_io_x3),
    .io_s(m_1243_io_s),
    .io_cout(m_1243_io_cout)
  );
  Adder m_1244 ( // @[MUL.scala 102:19]
    .io_x1(m_1244_io_x1),
    .io_x2(m_1244_io_x2),
    .io_x3(m_1244_io_x3),
    .io_s(m_1244_io_s),
    .io_cout(m_1244_io_cout)
  );
  Adder m_1245 ( // @[MUL.scala 102:19]
    .io_x1(m_1245_io_x1),
    .io_x2(m_1245_io_x2),
    .io_x3(m_1245_io_x3),
    .io_s(m_1245_io_s),
    .io_cout(m_1245_io_cout)
  );
  Adder m_1246 ( // @[MUL.scala 102:19]
    .io_x1(m_1246_io_x1),
    .io_x2(m_1246_io_x2),
    .io_x3(m_1246_io_x3),
    .io_s(m_1246_io_s),
    .io_cout(m_1246_io_cout)
  );
  Adder m_1247 ( // @[MUL.scala 102:19]
    .io_x1(m_1247_io_x1),
    .io_x2(m_1247_io_x2),
    .io_x3(m_1247_io_x3),
    .io_s(m_1247_io_s),
    .io_cout(m_1247_io_cout)
  );
  Adder m_1248 ( // @[MUL.scala 102:19]
    .io_x1(m_1248_io_x1),
    .io_x2(m_1248_io_x2),
    .io_x3(m_1248_io_x3),
    .io_s(m_1248_io_s),
    .io_cout(m_1248_io_cout)
  );
  Adder m_1249 ( // @[MUL.scala 102:19]
    .io_x1(m_1249_io_x1),
    .io_x2(m_1249_io_x2),
    .io_x3(m_1249_io_x3),
    .io_s(m_1249_io_s),
    .io_cout(m_1249_io_cout)
  );
  Adder m_1250 ( // @[MUL.scala 102:19]
    .io_x1(m_1250_io_x1),
    .io_x2(m_1250_io_x2),
    .io_x3(m_1250_io_x3),
    .io_s(m_1250_io_s),
    .io_cout(m_1250_io_cout)
  );
  Adder m_1251 ( // @[MUL.scala 102:19]
    .io_x1(m_1251_io_x1),
    .io_x2(m_1251_io_x2),
    .io_x3(m_1251_io_x3),
    .io_s(m_1251_io_s),
    .io_cout(m_1251_io_cout)
  );
  Adder m_1252 ( // @[MUL.scala 102:19]
    .io_x1(m_1252_io_x1),
    .io_x2(m_1252_io_x2),
    .io_x3(m_1252_io_x3),
    .io_s(m_1252_io_s),
    .io_cout(m_1252_io_cout)
  );
  Adder m_1253 ( // @[MUL.scala 102:19]
    .io_x1(m_1253_io_x1),
    .io_x2(m_1253_io_x2),
    .io_x3(m_1253_io_x3),
    .io_s(m_1253_io_s),
    .io_cout(m_1253_io_cout)
  );
  Adder m_1254 ( // @[MUL.scala 102:19]
    .io_x1(m_1254_io_x1),
    .io_x2(m_1254_io_x2),
    .io_x3(m_1254_io_x3),
    .io_s(m_1254_io_s),
    .io_cout(m_1254_io_cout)
  );
  Adder m_1255 ( // @[MUL.scala 102:19]
    .io_x1(m_1255_io_x1),
    .io_x2(m_1255_io_x2),
    .io_x3(m_1255_io_x3),
    .io_s(m_1255_io_s),
    .io_cout(m_1255_io_cout)
  );
  Adder m_1256 ( // @[MUL.scala 102:19]
    .io_x1(m_1256_io_x1),
    .io_x2(m_1256_io_x2),
    .io_x3(m_1256_io_x3),
    .io_s(m_1256_io_s),
    .io_cout(m_1256_io_cout)
  );
  Adder m_1257 ( // @[MUL.scala 102:19]
    .io_x1(m_1257_io_x1),
    .io_x2(m_1257_io_x2),
    .io_x3(m_1257_io_x3),
    .io_s(m_1257_io_s),
    .io_cout(m_1257_io_cout)
  );
  Adder m_1258 ( // @[MUL.scala 102:19]
    .io_x1(m_1258_io_x1),
    .io_x2(m_1258_io_x2),
    .io_x3(m_1258_io_x3),
    .io_s(m_1258_io_s),
    .io_cout(m_1258_io_cout)
  );
  Adder m_1259 ( // @[MUL.scala 102:19]
    .io_x1(m_1259_io_x1),
    .io_x2(m_1259_io_x2),
    .io_x3(m_1259_io_x3),
    .io_s(m_1259_io_s),
    .io_cout(m_1259_io_cout)
  );
  Adder m_1260 ( // @[MUL.scala 102:19]
    .io_x1(m_1260_io_x1),
    .io_x2(m_1260_io_x2),
    .io_x3(m_1260_io_x3),
    .io_s(m_1260_io_s),
    .io_cout(m_1260_io_cout)
  );
  Adder m_1261 ( // @[MUL.scala 102:19]
    .io_x1(m_1261_io_x1),
    .io_x2(m_1261_io_x2),
    .io_x3(m_1261_io_x3),
    .io_s(m_1261_io_s),
    .io_cout(m_1261_io_cout)
  );
  Adder m_1262 ( // @[MUL.scala 102:19]
    .io_x1(m_1262_io_x1),
    .io_x2(m_1262_io_x2),
    .io_x3(m_1262_io_x3),
    .io_s(m_1262_io_s),
    .io_cout(m_1262_io_cout)
  );
  Adder m_1263 ( // @[MUL.scala 102:19]
    .io_x1(m_1263_io_x1),
    .io_x2(m_1263_io_x2),
    .io_x3(m_1263_io_x3),
    .io_s(m_1263_io_s),
    .io_cout(m_1263_io_cout)
  );
  Adder m_1264 ( // @[MUL.scala 102:19]
    .io_x1(m_1264_io_x1),
    .io_x2(m_1264_io_x2),
    .io_x3(m_1264_io_x3),
    .io_s(m_1264_io_s),
    .io_cout(m_1264_io_cout)
  );
  Adder m_1265 ( // @[MUL.scala 102:19]
    .io_x1(m_1265_io_x1),
    .io_x2(m_1265_io_x2),
    .io_x3(m_1265_io_x3),
    .io_s(m_1265_io_s),
    .io_cout(m_1265_io_cout)
  );
  Adder m_1266 ( // @[MUL.scala 102:19]
    .io_x1(m_1266_io_x1),
    .io_x2(m_1266_io_x2),
    .io_x3(m_1266_io_x3),
    .io_s(m_1266_io_s),
    .io_cout(m_1266_io_cout)
  );
  Adder m_1267 ( // @[MUL.scala 102:19]
    .io_x1(m_1267_io_x1),
    .io_x2(m_1267_io_x2),
    .io_x3(m_1267_io_x3),
    .io_s(m_1267_io_s),
    .io_cout(m_1267_io_cout)
  );
  Adder m_1268 ( // @[MUL.scala 102:19]
    .io_x1(m_1268_io_x1),
    .io_x2(m_1268_io_x2),
    .io_x3(m_1268_io_x3),
    .io_s(m_1268_io_s),
    .io_cout(m_1268_io_cout)
  );
  Adder m_1269 ( // @[MUL.scala 102:19]
    .io_x1(m_1269_io_x1),
    .io_x2(m_1269_io_x2),
    .io_x3(m_1269_io_x3),
    .io_s(m_1269_io_s),
    .io_cout(m_1269_io_cout)
  );
  Half_Adder m_1270 ( // @[MUL.scala 124:19]
    .io_in_0(m_1270_io_in_0),
    .io_in_1(m_1270_io_in_1),
    .io_out_0(m_1270_io_out_0),
    .io_out_1(m_1270_io_out_1)
  );
  Adder m_1271 ( // @[MUL.scala 102:19]
    .io_x1(m_1271_io_x1),
    .io_x2(m_1271_io_x2),
    .io_x3(m_1271_io_x3),
    .io_s(m_1271_io_s),
    .io_cout(m_1271_io_cout)
  );
  Adder m_1272 ( // @[MUL.scala 102:19]
    .io_x1(m_1272_io_x1),
    .io_x2(m_1272_io_x2),
    .io_x3(m_1272_io_x3),
    .io_s(m_1272_io_s),
    .io_cout(m_1272_io_cout)
  );
  Adder m_1273 ( // @[MUL.scala 102:19]
    .io_x1(m_1273_io_x1),
    .io_x2(m_1273_io_x2),
    .io_x3(m_1273_io_x3),
    .io_s(m_1273_io_s),
    .io_cout(m_1273_io_cout)
  );
  Adder m_1274 ( // @[MUL.scala 102:19]
    .io_x1(m_1274_io_x1),
    .io_x2(m_1274_io_x2),
    .io_x3(m_1274_io_x3),
    .io_s(m_1274_io_s),
    .io_cout(m_1274_io_cout)
  );
  Adder m_1275 ( // @[MUL.scala 102:19]
    .io_x1(m_1275_io_x1),
    .io_x2(m_1275_io_x2),
    .io_x3(m_1275_io_x3),
    .io_s(m_1275_io_s),
    .io_cout(m_1275_io_cout)
  );
  Adder m_1276 ( // @[MUL.scala 102:19]
    .io_x1(m_1276_io_x1),
    .io_x2(m_1276_io_x2),
    .io_x3(m_1276_io_x3),
    .io_s(m_1276_io_s),
    .io_cout(m_1276_io_cout)
  );
  Adder m_1277 ( // @[MUL.scala 102:19]
    .io_x1(m_1277_io_x1),
    .io_x2(m_1277_io_x2),
    .io_x3(m_1277_io_x3),
    .io_s(m_1277_io_s),
    .io_cout(m_1277_io_cout)
  );
  Adder m_1278 ( // @[MUL.scala 102:19]
    .io_x1(m_1278_io_x1),
    .io_x2(m_1278_io_x2),
    .io_x3(m_1278_io_x3),
    .io_s(m_1278_io_s),
    .io_cout(m_1278_io_cout)
  );
  Adder m_1279 ( // @[MUL.scala 102:19]
    .io_x1(m_1279_io_x1),
    .io_x2(m_1279_io_x2),
    .io_x3(m_1279_io_x3),
    .io_s(m_1279_io_s),
    .io_cout(m_1279_io_cout)
  );
  Adder m_1280 ( // @[MUL.scala 102:19]
    .io_x1(m_1280_io_x1),
    .io_x2(m_1280_io_x2),
    .io_x3(m_1280_io_x3),
    .io_s(m_1280_io_s),
    .io_cout(m_1280_io_cout)
  );
  Adder m_1281 ( // @[MUL.scala 102:19]
    .io_x1(m_1281_io_x1),
    .io_x2(m_1281_io_x2),
    .io_x3(m_1281_io_x3),
    .io_s(m_1281_io_s),
    .io_cout(m_1281_io_cout)
  );
  Adder m_1282 ( // @[MUL.scala 102:19]
    .io_x1(m_1282_io_x1),
    .io_x2(m_1282_io_x2),
    .io_x3(m_1282_io_x3),
    .io_s(m_1282_io_s),
    .io_cout(m_1282_io_cout)
  );
  Adder m_1283 ( // @[MUL.scala 102:19]
    .io_x1(m_1283_io_x1),
    .io_x2(m_1283_io_x2),
    .io_x3(m_1283_io_x3),
    .io_s(m_1283_io_s),
    .io_cout(m_1283_io_cout)
  );
  Adder m_1284 ( // @[MUL.scala 102:19]
    .io_x1(m_1284_io_x1),
    .io_x2(m_1284_io_x2),
    .io_x3(m_1284_io_x3),
    .io_s(m_1284_io_s),
    .io_cout(m_1284_io_cout)
  );
  Adder m_1285 ( // @[MUL.scala 102:19]
    .io_x1(m_1285_io_x1),
    .io_x2(m_1285_io_x2),
    .io_x3(m_1285_io_x3),
    .io_s(m_1285_io_s),
    .io_cout(m_1285_io_cout)
  );
  Adder m_1286 ( // @[MUL.scala 102:19]
    .io_x1(m_1286_io_x1),
    .io_x2(m_1286_io_x2),
    .io_x3(m_1286_io_x3),
    .io_s(m_1286_io_s),
    .io_cout(m_1286_io_cout)
  );
  Adder m_1287 ( // @[MUL.scala 102:19]
    .io_x1(m_1287_io_x1),
    .io_x2(m_1287_io_x2),
    .io_x3(m_1287_io_x3),
    .io_s(m_1287_io_s),
    .io_cout(m_1287_io_cout)
  );
  Adder m_1288 ( // @[MUL.scala 102:19]
    .io_x1(m_1288_io_x1),
    .io_x2(m_1288_io_x2),
    .io_x3(m_1288_io_x3),
    .io_s(m_1288_io_s),
    .io_cout(m_1288_io_cout)
  );
  Adder m_1289 ( // @[MUL.scala 102:19]
    .io_x1(m_1289_io_x1),
    .io_x2(m_1289_io_x2),
    .io_x3(m_1289_io_x3),
    .io_s(m_1289_io_s),
    .io_cout(m_1289_io_cout)
  );
  Adder m_1290 ( // @[MUL.scala 102:19]
    .io_x1(m_1290_io_x1),
    .io_x2(m_1290_io_x2),
    .io_x3(m_1290_io_x3),
    .io_s(m_1290_io_s),
    .io_cout(m_1290_io_cout)
  );
  Half_Adder m_1291 ( // @[MUL.scala 124:19]
    .io_in_0(m_1291_io_in_0),
    .io_in_1(m_1291_io_in_1),
    .io_out_0(m_1291_io_out_0),
    .io_out_1(m_1291_io_out_1)
  );
  Adder m_1292 ( // @[MUL.scala 102:19]
    .io_x1(m_1292_io_x1),
    .io_x2(m_1292_io_x2),
    .io_x3(m_1292_io_x3),
    .io_s(m_1292_io_s),
    .io_cout(m_1292_io_cout)
  );
  Adder m_1293 ( // @[MUL.scala 102:19]
    .io_x1(m_1293_io_x1),
    .io_x2(m_1293_io_x2),
    .io_x3(m_1293_io_x3),
    .io_s(m_1293_io_s),
    .io_cout(m_1293_io_cout)
  );
  Half_Adder m_1294 ( // @[MUL.scala 124:19]
    .io_in_0(m_1294_io_in_0),
    .io_in_1(m_1294_io_in_1),
    .io_out_0(m_1294_io_out_0),
    .io_out_1(m_1294_io_out_1)
  );
  Adder m_1295 ( // @[MUL.scala 102:19]
    .io_x1(m_1295_io_x1),
    .io_x2(m_1295_io_x2),
    .io_x3(m_1295_io_x3),
    .io_s(m_1295_io_s),
    .io_cout(m_1295_io_cout)
  );
  Adder m_1296 ( // @[MUL.scala 102:19]
    .io_x1(m_1296_io_x1),
    .io_x2(m_1296_io_x2),
    .io_x3(m_1296_io_x3),
    .io_s(m_1296_io_s),
    .io_cout(m_1296_io_cout)
  );
  Half_Adder m_1297 ( // @[MUL.scala 124:19]
    .io_in_0(m_1297_io_in_0),
    .io_in_1(m_1297_io_in_1),
    .io_out_0(m_1297_io_out_0),
    .io_out_1(m_1297_io_out_1)
  );
  Adder m_1298 ( // @[MUL.scala 102:19]
    .io_x1(m_1298_io_x1),
    .io_x2(m_1298_io_x2),
    .io_x3(m_1298_io_x3),
    .io_s(m_1298_io_s),
    .io_cout(m_1298_io_cout)
  );
  Adder m_1299 ( // @[MUL.scala 102:19]
    .io_x1(m_1299_io_x1),
    .io_x2(m_1299_io_x2),
    .io_x3(m_1299_io_x3),
    .io_s(m_1299_io_s),
    .io_cout(m_1299_io_cout)
  );
  Half_Adder m_1300 ( // @[MUL.scala 124:19]
    .io_in_0(m_1300_io_in_0),
    .io_in_1(m_1300_io_in_1),
    .io_out_0(m_1300_io_out_0),
    .io_out_1(m_1300_io_out_1)
  );
  Adder m_1301 ( // @[MUL.scala 102:19]
    .io_x1(m_1301_io_x1),
    .io_x2(m_1301_io_x2),
    .io_x3(m_1301_io_x3),
    .io_s(m_1301_io_s),
    .io_cout(m_1301_io_cout)
  );
  Adder m_1302 ( // @[MUL.scala 102:19]
    .io_x1(m_1302_io_x1),
    .io_x2(m_1302_io_x2),
    .io_x3(m_1302_io_x3),
    .io_s(m_1302_io_s),
    .io_cout(m_1302_io_cout)
  );
  Half_Adder m_1303 ( // @[MUL.scala 124:19]
    .io_in_0(m_1303_io_in_0),
    .io_in_1(m_1303_io_in_1),
    .io_out_0(m_1303_io_out_0),
    .io_out_1(m_1303_io_out_1)
  );
  Adder m_1304 ( // @[MUL.scala 102:19]
    .io_x1(m_1304_io_x1),
    .io_x2(m_1304_io_x2),
    .io_x3(m_1304_io_x3),
    .io_s(m_1304_io_s),
    .io_cout(m_1304_io_cout)
  );
  Adder m_1305 ( // @[MUL.scala 102:19]
    .io_x1(m_1305_io_x1),
    .io_x2(m_1305_io_x2),
    .io_x3(m_1305_io_x3),
    .io_s(m_1305_io_s),
    .io_cout(m_1305_io_cout)
  );
  Adder m_1306 ( // @[MUL.scala 102:19]
    .io_x1(m_1306_io_x1),
    .io_x2(m_1306_io_x2),
    .io_x3(m_1306_io_x3),
    .io_s(m_1306_io_s),
    .io_cout(m_1306_io_cout)
  );
  Adder m_1307 ( // @[MUL.scala 102:19]
    .io_x1(m_1307_io_x1),
    .io_x2(m_1307_io_x2),
    .io_x3(m_1307_io_x3),
    .io_s(m_1307_io_s),
    .io_cout(m_1307_io_cout)
  );
  Adder m_1308 ( // @[MUL.scala 102:19]
    .io_x1(m_1308_io_x1),
    .io_x2(m_1308_io_x2),
    .io_x3(m_1308_io_x3),
    .io_s(m_1308_io_s),
    .io_cout(m_1308_io_cout)
  );
  Adder m_1309 ( // @[MUL.scala 102:19]
    .io_x1(m_1309_io_x1),
    .io_x2(m_1309_io_x2),
    .io_x3(m_1309_io_x3),
    .io_s(m_1309_io_s),
    .io_cout(m_1309_io_cout)
  );
  Adder m_1310 ( // @[MUL.scala 102:19]
    .io_x1(m_1310_io_x1),
    .io_x2(m_1310_io_x2),
    .io_x3(m_1310_io_x3),
    .io_s(m_1310_io_s),
    .io_cout(m_1310_io_cout)
  );
  Adder m_1311 ( // @[MUL.scala 102:19]
    .io_x1(m_1311_io_x1),
    .io_x2(m_1311_io_x2),
    .io_x3(m_1311_io_x3),
    .io_s(m_1311_io_s),
    .io_cout(m_1311_io_cout)
  );
  Adder m_1312 ( // @[MUL.scala 102:19]
    .io_x1(m_1312_io_x1),
    .io_x2(m_1312_io_x2),
    .io_x3(m_1312_io_x3),
    .io_s(m_1312_io_s),
    .io_cout(m_1312_io_cout)
  );
  Adder m_1313 ( // @[MUL.scala 102:19]
    .io_x1(m_1313_io_x1),
    .io_x2(m_1313_io_x2),
    .io_x3(m_1313_io_x3),
    .io_s(m_1313_io_s),
    .io_cout(m_1313_io_cout)
  );
  Adder m_1314 ( // @[MUL.scala 102:19]
    .io_x1(m_1314_io_x1),
    .io_x2(m_1314_io_x2),
    .io_x3(m_1314_io_x3),
    .io_s(m_1314_io_s),
    .io_cout(m_1314_io_cout)
  );
  Adder m_1315 ( // @[MUL.scala 102:19]
    .io_x1(m_1315_io_x1),
    .io_x2(m_1315_io_x2),
    .io_x3(m_1315_io_x3),
    .io_s(m_1315_io_s),
    .io_cout(m_1315_io_cout)
  );
  Adder m_1316 ( // @[MUL.scala 102:19]
    .io_x1(m_1316_io_x1),
    .io_x2(m_1316_io_x2),
    .io_x3(m_1316_io_x3),
    .io_s(m_1316_io_s),
    .io_cout(m_1316_io_cout)
  );
  Half_Adder m_1317 ( // @[MUL.scala 124:19]
    .io_in_0(m_1317_io_in_0),
    .io_in_1(m_1317_io_in_1),
    .io_out_0(m_1317_io_out_0),
    .io_out_1(m_1317_io_out_1)
  );
  Adder m_1318 ( // @[MUL.scala 102:19]
    .io_x1(m_1318_io_x1),
    .io_x2(m_1318_io_x2),
    .io_x3(m_1318_io_x3),
    .io_s(m_1318_io_s),
    .io_cout(m_1318_io_cout)
  );
  Adder m_1319 ( // @[MUL.scala 102:19]
    .io_x1(m_1319_io_x1),
    .io_x2(m_1319_io_x2),
    .io_x3(m_1319_io_x3),
    .io_s(m_1319_io_s),
    .io_cout(m_1319_io_cout)
  );
  Adder m_1320 ( // @[MUL.scala 102:19]
    .io_x1(m_1320_io_x1),
    .io_x2(m_1320_io_x2),
    .io_x3(m_1320_io_x3),
    .io_s(m_1320_io_s),
    .io_cout(m_1320_io_cout)
  );
  Adder m_1321 ( // @[MUL.scala 102:19]
    .io_x1(m_1321_io_x1),
    .io_x2(m_1321_io_x2),
    .io_x3(m_1321_io_x3),
    .io_s(m_1321_io_s),
    .io_cout(m_1321_io_cout)
  );
  Adder m_1322 ( // @[MUL.scala 102:19]
    .io_x1(m_1322_io_x1),
    .io_x2(m_1322_io_x2),
    .io_x3(m_1322_io_x3),
    .io_s(m_1322_io_s),
    .io_cout(m_1322_io_cout)
  );
  Adder m_1323 ( // @[MUL.scala 102:19]
    .io_x1(m_1323_io_x1),
    .io_x2(m_1323_io_x2),
    .io_x3(m_1323_io_x3),
    .io_s(m_1323_io_s),
    .io_cout(m_1323_io_cout)
  );
  Half_Adder m_1324 ( // @[MUL.scala 124:19]
    .io_in_0(m_1324_io_in_0),
    .io_in_1(m_1324_io_in_1),
    .io_out_0(m_1324_io_out_0),
    .io_out_1(m_1324_io_out_1)
  );
  Half_Adder m_1325 ( // @[MUL.scala 124:19]
    .io_in_0(m_1325_io_in_0),
    .io_in_1(m_1325_io_in_1),
    .io_out_0(m_1325_io_out_0),
    .io_out_1(m_1325_io_out_1)
  );
  Half_Adder m_1326 ( // @[MUL.scala 124:19]
    .io_in_0(m_1326_io_in_0),
    .io_in_1(m_1326_io_in_1),
    .io_out_0(m_1326_io_out_0),
    .io_out_1(m_1326_io_out_1)
  );
  Half_Adder m_1327 ( // @[MUL.scala 124:19]
    .io_in_0(m_1327_io_in_0),
    .io_in_1(m_1327_io_in_1),
    .io_out_0(m_1327_io_out_0),
    .io_out_1(m_1327_io_out_1)
  );
  Half_Adder m_1328 ( // @[MUL.scala 124:19]
    .io_in_0(m_1328_io_in_0),
    .io_in_1(m_1328_io_in_1),
    .io_out_0(m_1328_io_out_0),
    .io_out_1(m_1328_io_out_1)
  );
  Half_Adder m_1329 ( // @[MUL.scala 124:19]
    .io_in_0(m_1329_io_in_0),
    .io_in_1(m_1329_io_in_1),
    .io_out_0(m_1329_io_out_0),
    .io_out_1(m_1329_io_out_1)
  );
  Half_Adder m_1330 ( // @[MUL.scala 124:19]
    .io_in_0(m_1330_io_in_0),
    .io_in_1(m_1330_io_in_1),
    .io_out_0(m_1330_io_out_0),
    .io_out_1(m_1330_io_out_1)
  );
  Half_Adder m_1331 ( // @[MUL.scala 124:19]
    .io_in_0(m_1331_io_in_0),
    .io_in_1(m_1331_io_in_1),
    .io_out_0(m_1331_io_out_0),
    .io_out_1(m_1331_io_out_1)
  );
  Half_Adder m_1332 ( // @[MUL.scala 124:19]
    .io_in_0(m_1332_io_in_0),
    .io_in_1(m_1332_io_in_1),
    .io_out_0(m_1332_io_out_0),
    .io_out_1(m_1332_io_out_1)
  );
  Half_Adder m_1333 ( // @[MUL.scala 124:19]
    .io_in_0(m_1333_io_in_0),
    .io_in_1(m_1333_io_in_1),
    .io_out_0(m_1333_io_out_0),
    .io_out_1(m_1333_io_out_1)
  );
  Adder m_1334 ( // @[MUL.scala 102:19]
    .io_x1(m_1334_io_x1),
    .io_x2(m_1334_io_x2),
    .io_x3(m_1334_io_x3),
    .io_s(m_1334_io_s),
    .io_cout(m_1334_io_cout)
  );
  Adder m_1335 ( // @[MUL.scala 102:19]
    .io_x1(m_1335_io_x1),
    .io_x2(m_1335_io_x2),
    .io_x3(m_1335_io_x3),
    .io_s(m_1335_io_s),
    .io_cout(m_1335_io_cout)
  );
  Adder m_1336 ( // @[MUL.scala 102:19]
    .io_x1(m_1336_io_x1),
    .io_x2(m_1336_io_x2),
    .io_x3(m_1336_io_x3),
    .io_s(m_1336_io_s),
    .io_cout(m_1336_io_cout)
  );
  Adder m_1337 ( // @[MUL.scala 102:19]
    .io_x1(m_1337_io_x1),
    .io_x2(m_1337_io_x2),
    .io_x3(m_1337_io_x3),
    .io_s(m_1337_io_s),
    .io_cout(m_1337_io_cout)
  );
  Adder m_1338 ( // @[MUL.scala 102:19]
    .io_x1(m_1338_io_x1),
    .io_x2(m_1338_io_x2),
    .io_x3(m_1338_io_x3),
    .io_s(m_1338_io_s),
    .io_cout(m_1338_io_cout)
  );
  Adder m_1339 ( // @[MUL.scala 102:19]
    .io_x1(m_1339_io_x1),
    .io_x2(m_1339_io_x2),
    .io_x3(m_1339_io_x3),
    .io_s(m_1339_io_s),
    .io_cout(m_1339_io_cout)
  );
  Adder m_1340 ( // @[MUL.scala 102:19]
    .io_x1(m_1340_io_x1),
    .io_x2(m_1340_io_x2),
    .io_x3(m_1340_io_x3),
    .io_s(m_1340_io_s),
    .io_cout(m_1340_io_cout)
  );
  Adder m_1341 ( // @[MUL.scala 102:19]
    .io_x1(m_1341_io_x1),
    .io_x2(m_1341_io_x2),
    .io_x3(m_1341_io_x3),
    .io_s(m_1341_io_s),
    .io_cout(m_1341_io_cout)
  );
  Adder m_1342 ( // @[MUL.scala 102:19]
    .io_x1(m_1342_io_x1),
    .io_x2(m_1342_io_x2),
    .io_x3(m_1342_io_x3),
    .io_s(m_1342_io_s),
    .io_cout(m_1342_io_cout)
  );
  Adder m_1343 ( // @[MUL.scala 102:19]
    .io_x1(m_1343_io_x1),
    .io_x2(m_1343_io_x2),
    .io_x3(m_1343_io_x3),
    .io_s(m_1343_io_s),
    .io_cout(m_1343_io_cout)
  );
  Half_Adder m_1344 ( // @[MUL.scala 124:19]
    .io_in_0(m_1344_io_in_0),
    .io_in_1(m_1344_io_in_1),
    .io_out_0(m_1344_io_out_0),
    .io_out_1(m_1344_io_out_1)
  );
  Adder m_1345 ( // @[MUL.scala 102:19]
    .io_x1(m_1345_io_x1),
    .io_x2(m_1345_io_x2),
    .io_x3(m_1345_io_x3),
    .io_s(m_1345_io_s),
    .io_cout(m_1345_io_cout)
  );
  Half_Adder m_1346 ( // @[MUL.scala 124:19]
    .io_in_0(m_1346_io_in_0),
    .io_in_1(m_1346_io_in_1),
    .io_out_0(m_1346_io_out_0),
    .io_out_1(m_1346_io_out_1)
  );
  Adder m_1347 ( // @[MUL.scala 102:19]
    .io_x1(m_1347_io_x1),
    .io_x2(m_1347_io_x2),
    .io_x3(m_1347_io_x3),
    .io_s(m_1347_io_s),
    .io_cout(m_1347_io_cout)
  );
  Half_Adder m_1348 ( // @[MUL.scala 124:19]
    .io_in_0(m_1348_io_in_0),
    .io_in_1(m_1348_io_in_1),
    .io_out_0(m_1348_io_out_0),
    .io_out_1(m_1348_io_out_1)
  );
  Adder m_1349 ( // @[MUL.scala 102:19]
    .io_x1(m_1349_io_x1),
    .io_x2(m_1349_io_x2),
    .io_x3(m_1349_io_x3),
    .io_s(m_1349_io_s),
    .io_cout(m_1349_io_cout)
  );
  Half_Adder m_1350 ( // @[MUL.scala 124:19]
    .io_in_0(m_1350_io_in_0),
    .io_in_1(m_1350_io_in_1),
    .io_out_0(m_1350_io_out_0),
    .io_out_1(m_1350_io_out_1)
  );
  Adder m_1351 ( // @[MUL.scala 102:19]
    .io_x1(m_1351_io_x1),
    .io_x2(m_1351_io_x2),
    .io_x3(m_1351_io_x3),
    .io_s(m_1351_io_s),
    .io_cout(m_1351_io_cout)
  );
  Adder m_1352 ( // @[MUL.scala 102:19]
    .io_x1(m_1352_io_x1),
    .io_x2(m_1352_io_x2),
    .io_x3(m_1352_io_x3),
    .io_s(m_1352_io_s),
    .io_cout(m_1352_io_cout)
  );
  Adder m_1353 ( // @[MUL.scala 102:19]
    .io_x1(m_1353_io_x1),
    .io_x2(m_1353_io_x2),
    .io_x3(m_1353_io_x3),
    .io_s(m_1353_io_s),
    .io_cout(m_1353_io_cout)
  );
  Adder m_1354 ( // @[MUL.scala 102:19]
    .io_x1(m_1354_io_x1),
    .io_x2(m_1354_io_x2),
    .io_x3(m_1354_io_x3),
    .io_s(m_1354_io_s),
    .io_cout(m_1354_io_cout)
  );
  Adder m_1355 ( // @[MUL.scala 102:19]
    .io_x1(m_1355_io_x1),
    .io_x2(m_1355_io_x2),
    .io_x3(m_1355_io_x3),
    .io_s(m_1355_io_s),
    .io_cout(m_1355_io_cout)
  );
  Adder m_1356 ( // @[MUL.scala 102:19]
    .io_x1(m_1356_io_x1),
    .io_x2(m_1356_io_x2),
    .io_x3(m_1356_io_x3),
    .io_s(m_1356_io_s),
    .io_cout(m_1356_io_cout)
  );
  Adder m_1357 ( // @[MUL.scala 102:19]
    .io_x1(m_1357_io_x1),
    .io_x2(m_1357_io_x2),
    .io_x3(m_1357_io_x3),
    .io_s(m_1357_io_s),
    .io_cout(m_1357_io_cout)
  );
  Adder m_1358 ( // @[MUL.scala 102:19]
    .io_x1(m_1358_io_x1),
    .io_x2(m_1358_io_x2),
    .io_x3(m_1358_io_x3),
    .io_s(m_1358_io_s),
    .io_cout(m_1358_io_cout)
  );
  Adder m_1359 ( // @[MUL.scala 102:19]
    .io_x1(m_1359_io_x1),
    .io_x2(m_1359_io_x2),
    .io_x3(m_1359_io_x3),
    .io_s(m_1359_io_s),
    .io_cout(m_1359_io_cout)
  );
  Adder m_1360 ( // @[MUL.scala 102:19]
    .io_x1(m_1360_io_x1),
    .io_x2(m_1360_io_x2),
    .io_x3(m_1360_io_x3),
    .io_s(m_1360_io_s),
    .io_cout(m_1360_io_cout)
  );
  Adder m_1361 ( // @[MUL.scala 102:19]
    .io_x1(m_1361_io_x1),
    .io_x2(m_1361_io_x2),
    .io_x3(m_1361_io_x3),
    .io_s(m_1361_io_s),
    .io_cout(m_1361_io_cout)
  );
  Adder m_1362 ( // @[MUL.scala 102:19]
    .io_x1(m_1362_io_x1),
    .io_x2(m_1362_io_x2),
    .io_x3(m_1362_io_x3),
    .io_s(m_1362_io_s),
    .io_cout(m_1362_io_cout)
  );
  Adder m_1363 ( // @[MUL.scala 102:19]
    .io_x1(m_1363_io_x1),
    .io_x2(m_1363_io_x2),
    .io_x3(m_1363_io_x3),
    .io_s(m_1363_io_s),
    .io_cout(m_1363_io_cout)
  );
  Adder m_1364 ( // @[MUL.scala 102:19]
    .io_x1(m_1364_io_x1),
    .io_x2(m_1364_io_x2),
    .io_x3(m_1364_io_x3),
    .io_s(m_1364_io_s),
    .io_cout(m_1364_io_cout)
  );
  Adder m_1365 ( // @[MUL.scala 102:19]
    .io_x1(m_1365_io_x1),
    .io_x2(m_1365_io_x2),
    .io_x3(m_1365_io_x3),
    .io_s(m_1365_io_s),
    .io_cout(m_1365_io_cout)
  );
  Adder m_1366 ( // @[MUL.scala 102:19]
    .io_x1(m_1366_io_x1),
    .io_x2(m_1366_io_x2),
    .io_x3(m_1366_io_x3),
    .io_s(m_1366_io_s),
    .io_cout(m_1366_io_cout)
  );
  Adder m_1367 ( // @[MUL.scala 102:19]
    .io_x1(m_1367_io_x1),
    .io_x2(m_1367_io_x2),
    .io_x3(m_1367_io_x3),
    .io_s(m_1367_io_s),
    .io_cout(m_1367_io_cout)
  );
  Adder m_1368 ( // @[MUL.scala 102:19]
    .io_x1(m_1368_io_x1),
    .io_x2(m_1368_io_x2),
    .io_x3(m_1368_io_x3),
    .io_s(m_1368_io_s),
    .io_cout(m_1368_io_cout)
  );
  Adder m_1369 ( // @[MUL.scala 102:19]
    .io_x1(m_1369_io_x1),
    .io_x2(m_1369_io_x2),
    .io_x3(m_1369_io_x3),
    .io_s(m_1369_io_s),
    .io_cout(m_1369_io_cout)
  );
  Adder m_1370 ( // @[MUL.scala 102:19]
    .io_x1(m_1370_io_x1),
    .io_x2(m_1370_io_x2),
    .io_x3(m_1370_io_x3),
    .io_s(m_1370_io_s),
    .io_cout(m_1370_io_cout)
  );
  Half_Adder m_1371 ( // @[MUL.scala 124:19]
    .io_in_0(m_1371_io_in_0),
    .io_in_1(m_1371_io_in_1),
    .io_out_0(m_1371_io_out_0),
    .io_out_1(m_1371_io_out_1)
  );
  Adder m_1372 ( // @[MUL.scala 102:19]
    .io_x1(m_1372_io_x1),
    .io_x2(m_1372_io_x2),
    .io_x3(m_1372_io_x3),
    .io_s(m_1372_io_s),
    .io_cout(m_1372_io_cout)
  );
  Adder m_1373 ( // @[MUL.scala 102:19]
    .io_x1(m_1373_io_x1),
    .io_x2(m_1373_io_x2),
    .io_x3(m_1373_io_x3),
    .io_s(m_1373_io_s),
    .io_cout(m_1373_io_cout)
  );
  Half_Adder m_1374 ( // @[MUL.scala 124:19]
    .io_in_0(m_1374_io_in_0),
    .io_in_1(m_1374_io_in_1),
    .io_out_0(m_1374_io_out_0),
    .io_out_1(m_1374_io_out_1)
  );
  Adder m_1375 ( // @[MUL.scala 102:19]
    .io_x1(m_1375_io_x1),
    .io_x2(m_1375_io_x2),
    .io_x3(m_1375_io_x3),
    .io_s(m_1375_io_s),
    .io_cout(m_1375_io_cout)
  );
  Adder m_1376 ( // @[MUL.scala 102:19]
    .io_x1(m_1376_io_x1),
    .io_x2(m_1376_io_x2),
    .io_x3(m_1376_io_x3),
    .io_s(m_1376_io_s),
    .io_cout(m_1376_io_cout)
  );
  Half_Adder m_1377 ( // @[MUL.scala 124:19]
    .io_in_0(m_1377_io_in_0),
    .io_in_1(m_1377_io_in_1),
    .io_out_0(m_1377_io_out_0),
    .io_out_1(m_1377_io_out_1)
  );
  Adder m_1378 ( // @[MUL.scala 102:19]
    .io_x1(m_1378_io_x1),
    .io_x2(m_1378_io_x2),
    .io_x3(m_1378_io_x3),
    .io_s(m_1378_io_s),
    .io_cout(m_1378_io_cout)
  );
  Adder m_1379 ( // @[MUL.scala 102:19]
    .io_x1(m_1379_io_x1),
    .io_x2(m_1379_io_x2),
    .io_x3(m_1379_io_x3),
    .io_s(m_1379_io_s),
    .io_cout(m_1379_io_cout)
  );
  Half_Adder m_1380 ( // @[MUL.scala 124:19]
    .io_in_0(m_1380_io_in_0),
    .io_in_1(m_1380_io_in_1),
    .io_out_0(m_1380_io_out_0),
    .io_out_1(m_1380_io_out_1)
  );
  Adder m_1381 ( // @[MUL.scala 102:19]
    .io_x1(m_1381_io_x1),
    .io_x2(m_1381_io_x2),
    .io_x3(m_1381_io_x3),
    .io_s(m_1381_io_s),
    .io_cout(m_1381_io_cout)
  );
  Adder m_1382 ( // @[MUL.scala 102:19]
    .io_x1(m_1382_io_x1),
    .io_x2(m_1382_io_x2),
    .io_x3(m_1382_io_x3),
    .io_s(m_1382_io_s),
    .io_cout(m_1382_io_cout)
  );
  Half_Adder m_1383 ( // @[MUL.scala 124:19]
    .io_in_0(m_1383_io_in_0),
    .io_in_1(m_1383_io_in_1),
    .io_out_0(m_1383_io_out_0),
    .io_out_1(m_1383_io_out_1)
  );
  Adder m_1384 ( // @[MUL.scala 102:19]
    .io_x1(m_1384_io_x1),
    .io_x2(m_1384_io_x2),
    .io_x3(m_1384_io_x3),
    .io_s(m_1384_io_s),
    .io_cout(m_1384_io_cout)
  );
  Adder m_1385 ( // @[MUL.scala 102:19]
    .io_x1(m_1385_io_x1),
    .io_x2(m_1385_io_x2),
    .io_x3(m_1385_io_x3),
    .io_s(m_1385_io_s),
    .io_cout(m_1385_io_cout)
  );
  Adder m_1386 ( // @[MUL.scala 102:19]
    .io_x1(m_1386_io_x1),
    .io_x2(m_1386_io_x2),
    .io_x3(m_1386_io_x3),
    .io_s(m_1386_io_s),
    .io_cout(m_1386_io_cout)
  );
  Adder m_1387 ( // @[MUL.scala 102:19]
    .io_x1(m_1387_io_x1),
    .io_x2(m_1387_io_x2),
    .io_x3(m_1387_io_x3),
    .io_s(m_1387_io_s),
    .io_cout(m_1387_io_cout)
  );
  Adder m_1388 ( // @[MUL.scala 102:19]
    .io_x1(m_1388_io_x1),
    .io_x2(m_1388_io_x2),
    .io_x3(m_1388_io_x3),
    .io_s(m_1388_io_s),
    .io_cout(m_1388_io_cout)
  );
  Adder m_1389 ( // @[MUL.scala 102:19]
    .io_x1(m_1389_io_x1),
    .io_x2(m_1389_io_x2),
    .io_x3(m_1389_io_x3),
    .io_s(m_1389_io_s),
    .io_cout(m_1389_io_cout)
  );
  Adder m_1390 ( // @[MUL.scala 102:19]
    .io_x1(m_1390_io_x1),
    .io_x2(m_1390_io_x2),
    .io_x3(m_1390_io_x3),
    .io_s(m_1390_io_s),
    .io_cout(m_1390_io_cout)
  );
  Adder m_1391 ( // @[MUL.scala 102:19]
    .io_x1(m_1391_io_x1),
    .io_x2(m_1391_io_x2),
    .io_x3(m_1391_io_x3),
    .io_s(m_1391_io_s),
    .io_cout(m_1391_io_cout)
  );
  Adder m_1392 ( // @[MUL.scala 102:19]
    .io_x1(m_1392_io_x1),
    .io_x2(m_1392_io_x2),
    .io_x3(m_1392_io_x3),
    .io_s(m_1392_io_s),
    .io_cout(m_1392_io_cout)
  );
  Adder m_1393 ( // @[MUL.scala 102:19]
    .io_x1(m_1393_io_x1),
    .io_x2(m_1393_io_x2),
    .io_x3(m_1393_io_x3),
    .io_s(m_1393_io_s),
    .io_cout(m_1393_io_cout)
  );
  Adder m_1394 ( // @[MUL.scala 102:19]
    .io_x1(m_1394_io_x1),
    .io_x2(m_1394_io_x2),
    .io_x3(m_1394_io_x3),
    .io_s(m_1394_io_s),
    .io_cout(m_1394_io_cout)
  );
  Adder m_1395 ( // @[MUL.scala 102:19]
    .io_x1(m_1395_io_x1),
    .io_x2(m_1395_io_x2),
    .io_x3(m_1395_io_x3),
    .io_s(m_1395_io_s),
    .io_cout(m_1395_io_cout)
  );
  Adder m_1396 ( // @[MUL.scala 102:19]
    .io_x1(m_1396_io_x1),
    .io_x2(m_1396_io_x2),
    .io_x3(m_1396_io_x3),
    .io_s(m_1396_io_s),
    .io_cout(m_1396_io_cout)
  );
  Adder m_1397 ( // @[MUL.scala 102:19]
    .io_x1(m_1397_io_x1),
    .io_x2(m_1397_io_x2),
    .io_x3(m_1397_io_x3),
    .io_s(m_1397_io_s),
    .io_cout(m_1397_io_cout)
  );
  Adder m_1398 ( // @[MUL.scala 102:19]
    .io_x1(m_1398_io_x1),
    .io_x2(m_1398_io_x2),
    .io_x3(m_1398_io_x3),
    .io_s(m_1398_io_s),
    .io_cout(m_1398_io_cout)
  );
  Adder m_1399 ( // @[MUL.scala 102:19]
    .io_x1(m_1399_io_x1),
    .io_x2(m_1399_io_x2),
    .io_x3(m_1399_io_x3),
    .io_s(m_1399_io_s),
    .io_cout(m_1399_io_cout)
  );
  Adder m_1400 ( // @[MUL.scala 102:19]
    .io_x1(m_1400_io_x1),
    .io_x2(m_1400_io_x2),
    .io_x3(m_1400_io_x3),
    .io_s(m_1400_io_s),
    .io_cout(m_1400_io_cout)
  );
  Adder m_1401 ( // @[MUL.scala 102:19]
    .io_x1(m_1401_io_x1),
    .io_x2(m_1401_io_x2),
    .io_x3(m_1401_io_x3),
    .io_s(m_1401_io_s),
    .io_cout(m_1401_io_cout)
  );
  Adder m_1402 ( // @[MUL.scala 102:19]
    .io_x1(m_1402_io_x1),
    .io_x2(m_1402_io_x2),
    .io_x3(m_1402_io_x3),
    .io_s(m_1402_io_s),
    .io_cout(m_1402_io_cout)
  );
  Adder m_1403 ( // @[MUL.scala 102:19]
    .io_x1(m_1403_io_x1),
    .io_x2(m_1403_io_x2),
    .io_x3(m_1403_io_x3),
    .io_s(m_1403_io_s),
    .io_cout(m_1403_io_cout)
  );
  Adder m_1404 ( // @[MUL.scala 102:19]
    .io_x1(m_1404_io_x1),
    .io_x2(m_1404_io_x2),
    .io_x3(m_1404_io_x3),
    .io_s(m_1404_io_s),
    .io_cout(m_1404_io_cout)
  );
  Adder m_1405 ( // @[MUL.scala 102:19]
    .io_x1(m_1405_io_x1),
    .io_x2(m_1405_io_x2),
    .io_x3(m_1405_io_x3),
    .io_s(m_1405_io_s),
    .io_cout(m_1405_io_cout)
  );
  Adder m_1406 ( // @[MUL.scala 102:19]
    .io_x1(m_1406_io_x1),
    .io_x2(m_1406_io_x2),
    .io_x3(m_1406_io_x3),
    .io_s(m_1406_io_s),
    .io_cout(m_1406_io_cout)
  );
  Adder m_1407 ( // @[MUL.scala 102:19]
    .io_x1(m_1407_io_x1),
    .io_x2(m_1407_io_x2),
    .io_x3(m_1407_io_x3),
    .io_s(m_1407_io_s),
    .io_cout(m_1407_io_cout)
  );
  Adder m_1408 ( // @[MUL.scala 102:19]
    .io_x1(m_1408_io_x1),
    .io_x2(m_1408_io_x2),
    .io_x3(m_1408_io_x3),
    .io_s(m_1408_io_s),
    .io_cout(m_1408_io_cout)
  );
  Adder m_1409 ( // @[MUL.scala 102:19]
    .io_x1(m_1409_io_x1),
    .io_x2(m_1409_io_x2),
    .io_x3(m_1409_io_x3),
    .io_s(m_1409_io_s),
    .io_cout(m_1409_io_cout)
  );
  Adder m_1410 ( // @[MUL.scala 102:19]
    .io_x1(m_1410_io_x1),
    .io_x2(m_1410_io_x2),
    .io_x3(m_1410_io_x3),
    .io_s(m_1410_io_s),
    .io_cout(m_1410_io_cout)
  );
  Adder m_1411 ( // @[MUL.scala 102:19]
    .io_x1(m_1411_io_x1),
    .io_x2(m_1411_io_x2),
    .io_x3(m_1411_io_x3),
    .io_s(m_1411_io_s),
    .io_cout(m_1411_io_cout)
  );
  Adder m_1412 ( // @[MUL.scala 102:19]
    .io_x1(m_1412_io_x1),
    .io_x2(m_1412_io_x2),
    .io_x3(m_1412_io_x3),
    .io_s(m_1412_io_s),
    .io_cout(m_1412_io_cout)
  );
  Adder m_1413 ( // @[MUL.scala 102:19]
    .io_x1(m_1413_io_x1),
    .io_x2(m_1413_io_x2),
    .io_x3(m_1413_io_x3),
    .io_s(m_1413_io_s),
    .io_cout(m_1413_io_cout)
  );
  Half_Adder m_1414 ( // @[MUL.scala 124:19]
    .io_in_0(m_1414_io_in_0),
    .io_in_1(m_1414_io_in_1),
    .io_out_0(m_1414_io_out_0),
    .io_out_1(m_1414_io_out_1)
  );
  Adder m_1415 ( // @[MUL.scala 102:19]
    .io_x1(m_1415_io_x1),
    .io_x2(m_1415_io_x2),
    .io_x3(m_1415_io_x3),
    .io_s(m_1415_io_s),
    .io_cout(m_1415_io_cout)
  );
  Adder m_1416 ( // @[MUL.scala 102:19]
    .io_x1(m_1416_io_x1),
    .io_x2(m_1416_io_x2),
    .io_x3(m_1416_io_x3),
    .io_s(m_1416_io_s),
    .io_cout(m_1416_io_cout)
  );
  Adder m_1417 ( // @[MUL.scala 102:19]
    .io_x1(m_1417_io_x1),
    .io_x2(m_1417_io_x2),
    .io_x3(m_1417_io_x3),
    .io_s(m_1417_io_s),
    .io_cout(m_1417_io_cout)
  );
  Half_Adder m_1418 ( // @[MUL.scala 124:19]
    .io_in_0(m_1418_io_in_0),
    .io_in_1(m_1418_io_in_1),
    .io_out_0(m_1418_io_out_0),
    .io_out_1(m_1418_io_out_1)
  );
  Adder m_1419 ( // @[MUL.scala 102:19]
    .io_x1(m_1419_io_x1),
    .io_x2(m_1419_io_x2),
    .io_x3(m_1419_io_x3),
    .io_s(m_1419_io_s),
    .io_cout(m_1419_io_cout)
  );
  Adder m_1420 ( // @[MUL.scala 102:19]
    .io_x1(m_1420_io_x1),
    .io_x2(m_1420_io_x2),
    .io_x3(m_1420_io_x3),
    .io_s(m_1420_io_s),
    .io_cout(m_1420_io_cout)
  );
  Adder m_1421 ( // @[MUL.scala 102:19]
    .io_x1(m_1421_io_x1),
    .io_x2(m_1421_io_x2),
    .io_x3(m_1421_io_x3),
    .io_s(m_1421_io_s),
    .io_cout(m_1421_io_cout)
  );
  Half_Adder m_1422 ( // @[MUL.scala 124:19]
    .io_in_0(m_1422_io_in_0),
    .io_in_1(m_1422_io_in_1),
    .io_out_0(m_1422_io_out_0),
    .io_out_1(m_1422_io_out_1)
  );
  Adder m_1423 ( // @[MUL.scala 102:19]
    .io_x1(m_1423_io_x1),
    .io_x2(m_1423_io_x2),
    .io_x3(m_1423_io_x3),
    .io_s(m_1423_io_s),
    .io_cout(m_1423_io_cout)
  );
  Adder m_1424 ( // @[MUL.scala 102:19]
    .io_x1(m_1424_io_x1),
    .io_x2(m_1424_io_x2),
    .io_x3(m_1424_io_x3),
    .io_s(m_1424_io_s),
    .io_cout(m_1424_io_cout)
  );
  Adder m_1425 ( // @[MUL.scala 102:19]
    .io_x1(m_1425_io_x1),
    .io_x2(m_1425_io_x2),
    .io_x3(m_1425_io_x3),
    .io_s(m_1425_io_s),
    .io_cout(m_1425_io_cout)
  );
  Half_Adder m_1426 ( // @[MUL.scala 124:19]
    .io_in_0(m_1426_io_in_0),
    .io_in_1(m_1426_io_in_1),
    .io_out_0(m_1426_io_out_0),
    .io_out_1(m_1426_io_out_1)
  );
  Adder m_1427 ( // @[MUL.scala 102:19]
    .io_x1(m_1427_io_x1),
    .io_x2(m_1427_io_x2),
    .io_x3(m_1427_io_x3),
    .io_s(m_1427_io_s),
    .io_cout(m_1427_io_cout)
  );
  Adder m_1428 ( // @[MUL.scala 102:19]
    .io_x1(m_1428_io_x1),
    .io_x2(m_1428_io_x2),
    .io_x3(m_1428_io_x3),
    .io_s(m_1428_io_s),
    .io_cout(m_1428_io_cout)
  );
  Adder m_1429 ( // @[MUL.scala 102:19]
    .io_x1(m_1429_io_x1),
    .io_x2(m_1429_io_x2),
    .io_x3(m_1429_io_x3),
    .io_s(m_1429_io_s),
    .io_cout(m_1429_io_cout)
  );
  Adder m_1430 ( // @[MUL.scala 102:19]
    .io_x1(m_1430_io_x1),
    .io_x2(m_1430_io_x2),
    .io_x3(m_1430_io_x3),
    .io_s(m_1430_io_s),
    .io_cout(m_1430_io_cout)
  );
  Adder m_1431 ( // @[MUL.scala 102:19]
    .io_x1(m_1431_io_x1),
    .io_x2(m_1431_io_x2),
    .io_x3(m_1431_io_x3),
    .io_s(m_1431_io_s),
    .io_cout(m_1431_io_cout)
  );
  Adder m_1432 ( // @[MUL.scala 102:19]
    .io_x1(m_1432_io_x1),
    .io_x2(m_1432_io_x2),
    .io_x3(m_1432_io_x3),
    .io_s(m_1432_io_s),
    .io_cout(m_1432_io_cout)
  );
  Adder m_1433 ( // @[MUL.scala 102:19]
    .io_x1(m_1433_io_x1),
    .io_x2(m_1433_io_x2),
    .io_x3(m_1433_io_x3),
    .io_s(m_1433_io_s),
    .io_cout(m_1433_io_cout)
  );
  Adder m_1434 ( // @[MUL.scala 102:19]
    .io_x1(m_1434_io_x1),
    .io_x2(m_1434_io_x2),
    .io_x3(m_1434_io_x3),
    .io_s(m_1434_io_s),
    .io_cout(m_1434_io_cout)
  );
  Adder m_1435 ( // @[MUL.scala 102:19]
    .io_x1(m_1435_io_x1),
    .io_x2(m_1435_io_x2),
    .io_x3(m_1435_io_x3),
    .io_s(m_1435_io_s),
    .io_cout(m_1435_io_cout)
  );
  Adder m_1436 ( // @[MUL.scala 102:19]
    .io_x1(m_1436_io_x1),
    .io_x2(m_1436_io_x2),
    .io_x3(m_1436_io_x3),
    .io_s(m_1436_io_s),
    .io_cout(m_1436_io_cout)
  );
  Adder m_1437 ( // @[MUL.scala 102:19]
    .io_x1(m_1437_io_x1),
    .io_x2(m_1437_io_x2),
    .io_x3(m_1437_io_x3),
    .io_s(m_1437_io_s),
    .io_cout(m_1437_io_cout)
  );
  Adder m_1438 ( // @[MUL.scala 102:19]
    .io_x1(m_1438_io_x1),
    .io_x2(m_1438_io_x2),
    .io_x3(m_1438_io_x3),
    .io_s(m_1438_io_s),
    .io_cout(m_1438_io_cout)
  );
  Adder m_1439 ( // @[MUL.scala 102:19]
    .io_x1(m_1439_io_x1),
    .io_x2(m_1439_io_x2),
    .io_x3(m_1439_io_x3),
    .io_s(m_1439_io_s),
    .io_cout(m_1439_io_cout)
  );
  Adder m_1440 ( // @[MUL.scala 102:19]
    .io_x1(m_1440_io_x1),
    .io_x2(m_1440_io_x2),
    .io_x3(m_1440_io_x3),
    .io_s(m_1440_io_s),
    .io_cout(m_1440_io_cout)
  );
  Adder m_1441 ( // @[MUL.scala 102:19]
    .io_x1(m_1441_io_x1),
    .io_x2(m_1441_io_x2),
    .io_x3(m_1441_io_x3),
    .io_s(m_1441_io_s),
    .io_cout(m_1441_io_cout)
  );
  Adder m_1442 ( // @[MUL.scala 102:19]
    .io_x1(m_1442_io_x1),
    .io_x2(m_1442_io_x2),
    .io_x3(m_1442_io_x3),
    .io_s(m_1442_io_s),
    .io_cout(m_1442_io_cout)
  );
  Adder m_1443 ( // @[MUL.scala 102:19]
    .io_x1(m_1443_io_x1),
    .io_x2(m_1443_io_x2),
    .io_x3(m_1443_io_x3),
    .io_s(m_1443_io_s),
    .io_cout(m_1443_io_cout)
  );
  Adder m_1444 ( // @[MUL.scala 102:19]
    .io_x1(m_1444_io_x1),
    .io_x2(m_1444_io_x2),
    .io_x3(m_1444_io_x3),
    .io_s(m_1444_io_s),
    .io_cout(m_1444_io_cout)
  );
  Adder m_1445 ( // @[MUL.scala 102:19]
    .io_x1(m_1445_io_x1),
    .io_x2(m_1445_io_x2),
    .io_x3(m_1445_io_x3),
    .io_s(m_1445_io_s),
    .io_cout(m_1445_io_cout)
  );
  Adder m_1446 ( // @[MUL.scala 102:19]
    .io_x1(m_1446_io_x1),
    .io_x2(m_1446_io_x2),
    .io_x3(m_1446_io_x3),
    .io_s(m_1446_io_s),
    .io_cout(m_1446_io_cout)
  );
  Adder m_1447 ( // @[MUL.scala 102:19]
    .io_x1(m_1447_io_x1),
    .io_x2(m_1447_io_x2),
    .io_x3(m_1447_io_x3),
    .io_s(m_1447_io_s),
    .io_cout(m_1447_io_cout)
  );
  Adder m_1448 ( // @[MUL.scala 102:19]
    .io_x1(m_1448_io_x1),
    .io_x2(m_1448_io_x2),
    .io_x3(m_1448_io_x3),
    .io_s(m_1448_io_s),
    .io_cout(m_1448_io_cout)
  );
  Adder m_1449 ( // @[MUL.scala 102:19]
    .io_x1(m_1449_io_x1),
    .io_x2(m_1449_io_x2),
    .io_x3(m_1449_io_x3),
    .io_s(m_1449_io_s),
    .io_cout(m_1449_io_cout)
  );
  Adder m_1450 ( // @[MUL.scala 102:19]
    .io_x1(m_1450_io_x1),
    .io_x2(m_1450_io_x2),
    .io_x3(m_1450_io_x3),
    .io_s(m_1450_io_s),
    .io_cout(m_1450_io_cout)
  );
  Adder m_1451 ( // @[MUL.scala 102:19]
    .io_x1(m_1451_io_x1),
    .io_x2(m_1451_io_x2),
    .io_x3(m_1451_io_x3),
    .io_s(m_1451_io_s),
    .io_cout(m_1451_io_cout)
  );
  Adder m_1452 ( // @[MUL.scala 102:19]
    .io_x1(m_1452_io_x1),
    .io_x2(m_1452_io_x2),
    .io_x3(m_1452_io_x3),
    .io_s(m_1452_io_s),
    .io_cout(m_1452_io_cout)
  );
  Adder m_1453 ( // @[MUL.scala 102:19]
    .io_x1(m_1453_io_x1),
    .io_x2(m_1453_io_x2),
    .io_x3(m_1453_io_x3),
    .io_s(m_1453_io_s),
    .io_cout(m_1453_io_cout)
  );
  Adder m_1454 ( // @[MUL.scala 102:19]
    .io_x1(m_1454_io_x1),
    .io_x2(m_1454_io_x2),
    .io_x3(m_1454_io_x3),
    .io_s(m_1454_io_s),
    .io_cout(m_1454_io_cout)
  );
  Adder m_1455 ( // @[MUL.scala 102:19]
    .io_x1(m_1455_io_x1),
    .io_x2(m_1455_io_x2),
    .io_x3(m_1455_io_x3),
    .io_s(m_1455_io_s),
    .io_cout(m_1455_io_cout)
  );
  Adder m_1456 ( // @[MUL.scala 102:19]
    .io_x1(m_1456_io_x1),
    .io_x2(m_1456_io_x2),
    .io_x3(m_1456_io_x3),
    .io_s(m_1456_io_s),
    .io_cout(m_1456_io_cout)
  );
  Adder m_1457 ( // @[MUL.scala 102:19]
    .io_x1(m_1457_io_x1),
    .io_x2(m_1457_io_x2),
    .io_x3(m_1457_io_x3),
    .io_s(m_1457_io_s),
    .io_cout(m_1457_io_cout)
  );
  Adder m_1458 ( // @[MUL.scala 102:19]
    .io_x1(m_1458_io_x1),
    .io_x2(m_1458_io_x2),
    .io_x3(m_1458_io_x3),
    .io_s(m_1458_io_s),
    .io_cout(m_1458_io_cout)
  );
  Adder m_1459 ( // @[MUL.scala 102:19]
    .io_x1(m_1459_io_x1),
    .io_x2(m_1459_io_x2),
    .io_x3(m_1459_io_x3),
    .io_s(m_1459_io_s),
    .io_cout(m_1459_io_cout)
  );
  Adder m_1460 ( // @[MUL.scala 102:19]
    .io_x1(m_1460_io_x1),
    .io_x2(m_1460_io_x2),
    .io_x3(m_1460_io_x3),
    .io_s(m_1460_io_s),
    .io_cout(m_1460_io_cout)
  );
  Adder m_1461 ( // @[MUL.scala 102:19]
    .io_x1(m_1461_io_x1),
    .io_x2(m_1461_io_x2),
    .io_x3(m_1461_io_x3),
    .io_s(m_1461_io_s),
    .io_cout(m_1461_io_cout)
  );
  Adder m_1462 ( // @[MUL.scala 102:19]
    .io_x1(m_1462_io_x1),
    .io_x2(m_1462_io_x2),
    .io_x3(m_1462_io_x3),
    .io_s(m_1462_io_s),
    .io_cout(m_1462_io_cout)
  );
  Adder m_1463 ( // @[MUL.scala 102:19]
    .io_x1(m_1463_io_x1),
    .io_x2(m_1463_io_x2),
    .io_x3(m_1463_io_x3),
    .io_s(m_1463_io_s),
    .io_cout(m_1463_io_cout)
  );
  Adder m_1464 ( // @[MUL.scala 102:19]
    .io_x1(m_1464_io_x1),
    .io_x2(m_1464_io_x2),
    .io_x3(m_1464_io_x3),
    .io_s(m_1464_io_s),
    .io_cout(m_1464_io_cout)
  );
  Adder m_1465 ( // @[MUL.scala 102:19]
    .io_x1(m_1465_io_x1),
    .io_x2(m_1465_io_x2),
    .io_x3(m_1465_io_x3),
    .io_s(m_1465_io_s),
    .io_cout(m_1465_io_cout)
  );
  Adder m_1466 ( // @[MUL.scala 102:19]
    .io_x1(m_1466_io_x1),
    .io_x2(m_1466_io_x2),
    .io_x3(m_1466_io_x3),
    .io_s(m_1466_io_s),
    .io_cout(m_1466_io_cout)
  );
  Half_Adder m_1467 ( // @[MUL.scala 124:19]
    .io_in_0(m_1467_io_in_0),
    .io_in_1(m_1467_io_in_1),
    .io_out_0(m_1467_io_out_0),
    .io_out_1(m_1467_io_out_1)
  );
  Adder m_1468 ( // @[MUL.scala 102:19]
    .io_x1(m_1468_io_x1),
    .io_x2(m_1468_io_x2),
    .io_x3(m_1468_io_x3),
    .io_s(m_1468_io_s),
    .io_cout(m_1468_io_cout)
  );
  Adder m_1469 ( // @[MUL.scala 102:19]
    .io_x1(m_1469_io_x1),
    .io_x2(m_1469_io_x2),
    .io_x3(m_1469_io_x3),
    .io_s(m_1469_io_s),
    .io_cout(m_1469_io_cout)
  );
  Adder m_1470 ( // @[MUL.scala 102:19]
    .io_x1(m_1470_io_x1),
    .io_x2(m_1470_io_x2),
    .io_x3(m_1470_io_x3),
    .io_s(m_1470_io_s),
    .io_cout(m_1470_io_cout)
  );
  Adder m_1471 ( // @[MUL.scala 102:19]
    .io_x1(m_1471_io_x1),
    .io_x2(m_1471_io_x2),
    .io_x3(m_1471_io_x3),
    .io_s(m_1471_io_s),
    .io_cout(m_1471_io_cout)
  );
  Half_Adder m_1472 ( // @[MUL.scala 124:19]
    .io_in_0(m_1472_io_in_0),
    .io_in_1(m_1472_io_in_1),
    .io_out_0(m_1472_io_out_0),
    .io_out_1(m_1472_io_out_1)
  );
  Adder m_1473 ( // @[MUL.scala 102:19]
    .io_x1(m_1473_io_x1),
    .io_x2(m_1473_io_x2),
    .io_x3(m_1473_io_x3),
    .io_s(m_1473_io_s),
    .io_cout(m_1473_io_cout)
  );
  Adder m_1474 ( // @[MUL.scala 102:19]
    .io_x1(m_1474_io_x1),
    .io_x2(m_1474_io_x2),
    .io_x3(m_1474_io_x3),
    .io_s(m_1474_io_s),
    .io_cout(m_1474_io_cout)
  );
  Adder m_1475 ( // @[MUL.scala 102:19]
    .io_x1(m_1475_io_x1),
    .io_x2(m_1475_io_x2),
    .io_x3(m_1475_io_x3),
    .io_s(m_1475_io_s),
    .io_cout(m_1475_io_cout)
  );
  Adder m_1476 ( // @[MUL.scala 102:19]
    .io_x1(m_1476_io_x1),
    .io_x2(m_1476_io_x2),
    .io_x3(m_1476_io_x3),
    .io_s(m_1476_io_s),
    .io_cout(m_1476_io_cout)
  );
  Half_Adder m_1477 ( // @[MUL.scala 124:19]
    .io_in_0(m_1477_io_in_0),
    .io_in_1(m_1477_io_in_1),
    .io_out_0(m_1477_io_out_0),
    .io_out_1(m_1477_io_out_1)
  );
  Adder m_1478 ( // @[MUL.scala 102:19]
    .io_x1(m_1478_io_x1),
    .io_x2(m_1478_io_x2),
    .io_x3(m_1478_io_x3),
    .io_s(m_1478_io_s),
    .io_cout(m_1478_io_cout)
  );
  Adder m_1479 ( // @[MUL.scala 102:19]
    .io_x1(m_1479_io_x1),
    .io_x2(m_1479_io_x2),
    .io_x3(m_1479_io_x3),
    .io_s(m_1479_io_s),
    .io_cout(m_1479_io_cout)
  );
  Adder m_1480 ( // @[MUL.scala 102:19]
    .io_x1(m_1480_io_x1),
    .io_x2(m_1480_io_x2),
    .io_x3(m_1480_io_x3),
    .io_s(m_1480_io_s),
    .io_cout(m_1480_io_cout)
  );
  Adder m_1481 ( // @[MUL.scala 102:19]
    .io_x1(m_1481_io_x1),
    .io_x2(m_1481_io_x2),
    .io_x3(m_1481_io_x3),
    .io_s(m_1481_io_s),
    .io_cout(m_1481_io_cout)
  );
  Half_Adder m_1482 ( // @[MUL.scala 124:19]
    .io_in_0(m_1482_io_in_0),
    .io_in_1(m_1482_io_in_1),
    .io_out_0(m_1482_io_out_0),
    .io_out_1(m_1482_io_out_1)
  );
  Adder m_1483 ( // @[MUL.scala 102:19]
    .io_x1(m_1483_io_x1),
    .io_x2(m_1483_io_x2),
    .io_x3(m_1483_io_x3),
    .io_s(m_1483_io_s),
    .io_cout(m_1483_io_cout)
  );
  Adder m_1484 ( // @[MUL.scala 102:19]
    .io_x1(m_1484_io_x1),
    .io_x2(m_1484_io_x2),
    .io_x3(m_1484_io_x3),
    .io_s(m_1484_io_s),
    .io_cout(m_1484_io_cout)
  );
  Adder m_1485 ( // @[MUL.scala 102:19]
    .io_x1(m_1485_io_x1),
    .io_x2(m_1485_io_x2),
    .io_x3(m_1485_io_x3),
    .io_s(m_1485_io_s),
    .io_cout(m_1485_io_cout)
  );
  Adder m_1486 ( // @[MUL.scala 102:19]
    .io_x1(m_1486_io_x1),
    .io_x2(m_1486_io_x2),
    .io_x3(m_1486_io_x3),
    .io_s(m_1486_io_s),
    .io_cout(m_1486_io_cout)
  );
  Half_Adder m_1487 ( // @[MUL.scala 124:19]
    .io_in_0(m_1487_io_in_0),
    .io_in_1(m_1487_io_in_1),
    .io_out_0(m_1487_io_out_0),
    .io_out_1(m_1487_io_out_1)
  );
  Adder m_1488 ( // @[MUL.scala 102:19]
    .io_x1(m_1488_io_x1),
    .io_x2(m_1488_io_x2),
    .io_x3(m_1488_io_x3),
    .io_s(m_1488_io_s),
    .io_cout(m_1488_io_cout)
  );
  Adder m_1489 ( // @[MUL.scala 102:19]
    .io_x1(m_1489_io_x1),
    .io_x2(m_1489_io_x2),
    .io_x3(m_1489_io_x3),
    .io_s(m_1489_io_s),
    .io_cout(m_1489_io_cout)
  );
  Adder m_1490 ( // @[MUL.scala 102:19]
    .io_x1(m_1490_io_x1),
    .io_x2(m_1490_io_x2),
    .io_x3(m_1490_io_x3),
    .io_s(m_1490_io_s),
    .io_cout(m_1490_io_cout)
  );
  Adder m_1491 ( // @[MUL.scala 102:19]
    .io_x1(m_1491_io_x1),
    .io_x2(m_1491_io_x2),
    .io_x3(m_1491_io_x3),
    .io_s(m_1491_io_s),
    .io_cout(m_1491_io_cout)
  );
  Adder m_1492 ( // @[MUL.scala 102:19]
    .io_x1(m_1492_io_x1),
    .io_x2(m_1492_io_x2),
    .io_x3(m_1492_io_x3),
    .io_s(m_1492_io_s),
    .io_cout(m_1492_io_cout)
  );
  Adder m_1493 ( // @[MUL.scala 102:19]
    .io_x1(m_1493_io_x1),
    .io_x2(m_1493_io_x2),
    .io_x3(m_1493_io_x3),
    .io_s(m_1493_io_s),
    .io_cout(m_1493_io_cout)
  );
  Adder m_1494 ( // @[MUL.scala 102:19]
    .io_x1(m_1494_io_x1),
    .io_x2(m_1494_io_x2),
    .io_x3(m_1494_io_x3),
    .io_s(m_1494_io_s),
    .io_cout(m_1494_io_cout)
  );
  Adder m_1495 ( // @[MUL.scala 102:19]
    .io_x1(m_1495_io_x1),
    .io_x2(m_1495_io_x2),
    .io_x3(m_1495_io_x3),
    .io_s(m_1495_io_s),
    .io_cout(m_1495_io_cout)
  );
  Adder m_1496 ( // @[MUL.scala 102:19]
    .io_x1(m_1496_io_x1),
    .io_x2(m_1496_io_x2),
    .io_x3(m_1496_io_x3),
    .io_s(m_1496_io_s),
    .io_cout(m_1496_io_cout)
  );
  Adder m_1497 ( // @[MUL.scala 102:19]
    .io_x1(m_1497_io_x1),
    .io_x2(m_1497_io_x2),
    .io_x3(m_1497_io_x3),
    .io_s(m_1497_io_s),
    .io_cout(m_1497_io_cout)
  );
  Adder m_1498 ( // @[MUL.scala 102:19]
    .io_x1(m_1498_io_x1),
    .io_x2(m_1498_io_x2),
    .io_x3(m_1498_io_x3),
    .io_s(m_1498_io_s),
    .io_cout(m_1498_io_cout)
  );
  Adder m_1499 ( // @[MUL.scala 102:19]
    .io_x1(m_1499_io_x1),
    .io_x2(m_1499_io_x2),
    .io_x3(m_1499_io_x3),
    .io_s(m_1499_io_s),
    .io_cout(m_1499_io_cout)
  );
  Adder m_1500 ( // @[MUL.scala 102:19]
    .io_x1(m_1500_io_x1),
    .io_x2(m_1500_io_x2),
    .io_x3(m_1500_io_x3),
    .io_s(m_1500_io_s),
    .io_cout(m_1500_io_cout)
  );
  Adder m_1501 ( // @[MUL.scala 102:19]
    .io_x1(m_1501_io_x1),
    .io_x2(m_1501_io_x2),
    .io_x3(m_1501_io_x3),
    .io_s(m_1501_io_s),
    .io_cout(m_1501_io_cout)
  );
  Adder m_1502 ( // @[MUL.scala 102:19]
    .io_x1(m_1502_io_x1),
    .io_x2(m_1502_io_x2),
    .io_x3(m_1502_io_x3),
    .io_s(m_1502_io_s),
    .io_cout(m_1502_io_cout)
  );
  Adder m_1503 ( // @[MUL.scala 102:19]
    .io_x1(m_1503_io_x1),
    .io_x2(m_1503_io_x2),
    .io_x3(m_1503_io_x3),
    .io_s(m_1503_io_s),
    .io_cout(m_1503_io_cout)
  );
  Adder m_1504 ( // @[MUL.scala 102:19]
    .io_x1(m_1504_io_x1),
    .io_x2(m_1504_io_x2),
    .io_x3(m_1504_io_x3),
    .io_s(m_1504_io_s),
    .io_cout(m_1504_io_cout)
  );
  Adder m_1505 ( // @[MUL.scala 102:19]
    .io_x1(m_1505_io_x1),
    .io_x2(m_1505_io_x2),
    .io_x3(m_1505_io_x3),
    .io_s(m_1505_io_s),
    .io_cout(m_1505_io_cout)
  );
  Adder m_1506 ( // @[MUL.scala 102:19]
    .io_x1(m_1506_io_x1),
    .io_x2(m_1506_io_x2),
    .io_x3(m_1506_io_x3),
    .io_s(m_1506_io_s),
    .io_cout(m_1506_io_cout)
  );
  Adder m_1507 ( // @[MUL.scala 102:19]
    .io_x1(m_1507_io_x1),
    .io_x2(m_1507_io_x2),
    .io_x3(m_1507_io_x3),
    .io_s(m_1507_io_s),
    .io_cout(m_1507_io_cout)
  );
  Adder m_1508 ( // @[MUL.scala 102:19]
    .io_x1(m_1508_io_x1),
    .io_x2(m_1508_io_x2),
    .io_x3(m_1508_io_x3),
    .io_s(m_1508_io_s),
    .io_cout(m_1508_io_cout)
  );
  Adder m_1509 ( // @[MUL.scala 102:19]
    .io_x1(m_1509_io_x1),
    .io_x2(m_1509_io_x2),
    .io_x3(m_1509_io_x3),
    .io_s(m_1509_io_s),
    .io_cout(m_1509_io_cout)
  );
  Adder m_1510 ( // @[MUL.scala 102:19]
    .io_x1(m_1510_io_x1),
    .io_x2(m_1510_io_x2),
    .io_x3(m_1510_io_x3),
    .io_s(m_1510_io_s),
    .io_cout(m_1510_io_cout)
  );
  Adder m_1511 ( // @[MUL.scala 102:19]
    .io_x1(m_1511_io_x1),
    .io_x2(m_1511_io_x2),
    .io_x3(m_1511_io_x3),
    .io_s(m_1511_io_s),
    .io_cout(m_1511_io_cout)
  );
  Adder m_1512 ( // @[MUL.scala 102:19]
    .io_x1(m_1512_io_x1),
    .io_x2(m_1512_io_x2),
    .io_x3(m_1512_io_x3),
    .io_s(m_1512_io_s),
    .io_cout(m_1512_io_cout)
  );
  Adder m_1513 ( // @[MUL.scala 102:19]
    .io_x1(m_1513_io_x1),
    .io_x2(m_1513_io_x2),
    .io_x3(m_1513_io_x3),
    .io_s(m_1513_io_s),
    .io_cout(m_1513_io_cout)
  );
  Adder m_1514 ( // @[MUL.scala 102:19]
    .io_x1(m_1514_io_x1),
    .io_x2(m_1514_io_x2),
    .io_x3(m_1514_io_x3),
    .io_s(m_1514_io_s),
    .io_cout(m_1514_io_cout)
  );
  Adder m_1515 ( // @[MUL.scala 102:19]
    .io_x1(m_1515_io_x1),
    .io_x2(m_1515_io_x2),
    .io_x3(m_1515_io_x3),
    .io_s(m_1515_io_s),
    .io_cout(m_1515_io_cout)
  );
  Adder m_1516 ( // @[MUL.scala 102:19]
    .io_x1(m_1516_io_x1),
    .io_x2(m_1516_io_x2),
    .io_x3(m_1516_io_x3),
    .io_s(m_1516_io_s),
    .io_cout(m_1516_io_cout)
  );
  Adder m_1517 ( // @[MUL.scala 102:19]
    .io_x1(m_1517_io_x1),
    .io_x2(m_1517_io_x2),
    .io_x3(m_1517_io_x3),
    .io_s(m_1517_io_s),
    .io_cout(m_1517_io_cout)
  );
  Adder m_1518 ( // @[MUL.scala 102:19]
    .io_x1(m_1518_io_x1),
    .io_x2(m_1518_io_x2),
    .io_x3(m_1518_io_x3),
    .io_s(m_1518_io_s),
    .io_cout(m_1518_io_cout)
  );
  Adder m_1519 ( // @[MUL.scala 102:19]
    .io_x1(m_1519_io_x1),
    .io_x2(m_1519_io_x2),
    .io_x3(m_1519_io_x3),
    .io_s(m_1519_io_s),
    .io_cout(m_1519_io_cout)
  );
  Adder m_1520 ( // @[MUL.scala 102:19]
    .io_x1(m_1520_io_x1),
    .io_x2(m_1520_io_x2),
    .io_x3(m_1520_io_x3),
    .io_s(m_1520_io_s),
    .io_cout(m_1520_io_cout)
  );
  Adder m_1521 ( // @[MUL.scala 102:19]
    .io_x1(m_1521_io_x1),
    .io_x2(m_1521_io_x2),
    .io_x3(m_1521_io_x3),
    .io_s(m_1521_io_s),
    .io_cout(m_1521_io_cout)
  );
  Adder m_1522 ( // @[MUL.scala 102:19]
    .io_x1(m_1522_io_x1),
    .io_x2(m_1522_io_x2),
    .io_x3(m_1522_io_x3),
    .io_s(m_1522_io_s),
    .io_cout(m_1522_io_cout)
  );
  Adder m_1523 ( // @[MUL.scala 102:19]
    .io_x1(m_1523_io_x1),
    .io_x2(m_1523_io_x2),
    .io_x3(m_1523_io_x3),
    .io_s(m_1523_io_s),
    .io_cout(m_1523_io_cout)
  );
  Adder m_1524 ( // @[MUL.scala 102:19]
    .io_x1(m_1524_io_x1),
    .io_x2(m_1524_io_x2),
    .io_x3(m_1524_io_x3),
    .io_s(m_1524_io_s),
    .io_cout(m_1524_io_cout)
  );
  Adder m_1525 ( // @[MUL.scala 102:19]
    .io_x1(m_1525_io_x1),
    .io_x2(m_1525_io_x2),
    .io_x3(m_1525_io_x3),
    .io_s(m_1525_io_s),
    .io_cout(m_1525_io_cout)
  );
  Adder m_1526 ( // @[MUL.scala 102:19]
    .io_x1(m_1526_io_x1),
    .io_x2(m_1526_io_x2),
    .io_x3(m_1526_io_x3),
    .io_s(m_1526_io_s),
    .io_cout(m_1526_io_cout)
  );
  Adder m_1527 ( // @[MUL.scala 102:19]
    .io_x1(m_1527_io_x1),
    .io_x2(m_1527_io_x2),
    .io_x3(m_1527_io_x3),
    .io_s(m_1527_io_s),
    .io_cout(m_1527_io_cout)
  );
  Adder m_1528 ( // @[MUL.scala 102:19]
    .io_x1(m_1528_io_x1),
    .io_x2(m_1528_io_x2),
    .io_x3(m_1528_io_x3),
    .io_s(m_1528_io_s),
    .io_cout(m_1528_io_cout)
  );
  Adder m_1529 ( // @[MUL.scala 102:19]
    .io_x1(m_1529_io_x1),
    .io_x2(m_1529_io_x2),
    .io_x3(m_1529_io_x3),
    .io_s(m_1529_io_s),
    .io_cout(m_1529_io_cout)
  );
  Adder m_1530 ( // @[MUL.scala 102:19]
    .io_x1(m_1530_io_x1),
    .io_x2(m_1530_io_x2),
    .io_x3(m_1530_io_x3),
    .io_s(m_1530_io_s),
    .io_cout(m_1530_io_cout)
  );
  Adder m_1531 ( // @[MUL.scala 102:19]
    .io_x1(m_1531_io_x1),
    .io_x2(m_1531_io_x2),
    .io_x3(m_1531_io_x3),
    .io_s(m_1531_io_s),
    .io_cout(m_1531_io_cout)
  );
  Adder m_1532 ( // @[MUL.scala 102:19]
    .io_x1(m_1532_io_x1),
    .io_x2(m_1532_io_x2),
    .io_x3(m_1532_io_x3),
    .io_s(m_1532_io_s),
    .io_cout(m_1532_io_cout)
  );
  Adder m_1533 ( // @[MUL.scala 102:19]
    .io_x1(m_1533_io_x1),
    .io_x2(m_1533_io_x2),
    .io_x3(m_1533_io_x3),
    .io_s(m_1533_io_s),
    .io_cout(m_1533_io_cout)
  );
  Adder m_1534 ( // @[MUL.scala 102:19]
    .io_x1(m_1534_io_x1),
    .io_x2(m_1534_io_x2),
    .io_x3(m_1534_io_x3),
    .io_s(m_1534_io_s),
    .io_cout(m_1534_io_cout)
  );
  Adder m_1535 ( // @[MUL.scala 102:19]
    .io_x1(m_1535_io_x1),
    .io_x2(m_1535_io_x2),
    .io_x3(m_1535_io_x3),
    .io_s(m_1535_io_s),
    .io_cout(m_1535_io_cout)
  );
  Adder m_1536 ( // @[MUL.scala 102:19]
    .io_x1(m_1536_io_x1),
    .io_x2(m_1536_io_x2),
    .io_x3(m_1536_io_x3),
    .io_s(m_1536_io_s),
    .io_cout(m_1536_io_cout)
  );
  Adder m_1537 ( // @[MUL.scala 102:19]
    .io_x1(m_1537_io_x1),
    .io_x2(m_1537_io_x2),
    .io_x3(m_1537_io_x3),
    .io_s(m_1537_io_s),
    .io_cout(m_1537_io_cout)
  );
  Adder m_1538 ( // @[MUL.scala 102:19]
    .io_x1(m_1538_io_x1),
    .io_x2(m_1538_io_x2),
    .io_x3(m_1538_io_x3),
    .io_s(m_1538_io_s),
    .io_cout(m_1538_io_cout)
  );
  Adder m_1539 ( // @[MUL.scala 102:19]
    .io_x1(m_1539_io_x1),
    .io_x2(m_1539_io_x2),
    .io_x3(m_1539_io_x3),
    .io_s(m_1539_io_s),
    .io_cout(m_1539_io_cout)
  );
  Adder m_1540 ( // @[MUL.scala 102:19]
    .io_x1(m_1540_io_x1),
    .io_x2(m_1540_io_x2),
    .io_x3(m_1540_io_x3),
    .io_s(m_1540_io_s),
    .io_cout(m_1540_io_cout)
  );
  Adder m_1541 ( // @[MUL.scala 102:19]
    .io_x1(m_1541_io_x1),
    .io_x2(m_1541_io_x2),
    .io_x3(m_1541_io_x3),
    .io_s(m_1541_io_s),
    .io_cout(m_1541_io_cout)
  );
  Half_Adder m_1542 ( // @[MUL.scala 124:19]
    .io_in_0(m_1542_io_in_0),
    .io_in_1(m_1542_io_in_1),
    .io_out_0(m_1542_io_out_0),
    .io_out_1(m_1542_io_out_1)
  );
  Adder m_1543 ( // @[MUL.scala 102:19]
    .io_x1(m_1543_io_x1),
    .io_x2(m_1543_io_x2),
    .io_x3(m_1543_io_x3),
    .io_s(m_1543_io_s),
    .io_cout(m_1543_io_cout)
  );
  Adder m_1544 ( // @[MUL.scala 102:19]
    .io_x1(m_1544_io_x1),
    .io_x2(m_1544_io_x2),
    .io_x3(m_1544_io_x3),
    .io_s(m_1544_io_s),
    .io_cout(m_1544_io_cout)
  );
  Adder m_1545 ( // @[MUL.scala 102:19]
    .io_x1(m_1545_io_x1),
    .io_x2(m_1545_io_x2),
    .io_x3(m_1545_io_x3),
    .io_s(m_1545_io_s),
    .io_cout(m_1545_io_cout)
  );
  Adder m_1546 ( // @[MUL.scala 102:19]
    .io_x1(m_1546_io_x1),
    .io_x2(m_1546_io_x2),
    .io_x3(m_1546_io_x3),
    .io_s(m_1546_io_s),
    .io_cout(m_1546_io_cout)
  );
  Half_Adder m_1547 ( // @[MUL.scala 124:19]
    .io_in_0(m_1547_io_in_0),
    .io_in_1(m_1547_io_in_1),
    .io_out_0(m_1547_io_out_0),
    .io_out_1(m_1547_io_out_1)
  );
  Adder m_1548 ( // @[MUL.scala 102:19]
    .io_x1(m_1548_io_x1),
    .io_x2(m_1548_io_x2),
    .io_x3(m_1548_io_x3),
    .io_s(m_1548_io_s),
    .io_cout(m_1548_io_cout)
  );
  Adder m_1549 ( // @[MUL.scala 102:19]
    .io_x1(m_1549_io_x1),
    .io_x2(m_1549_io_x2),
    .io_x3(m_1549_io_x3),
    .io_s(m_1549_io_s),
    .io_cout(m_1549_io_cout)
  );
  Adder m_1550 ( // @[MUL.scala 102:19]
    .io_x1(m_1550_io_x1),
    .io_x2(m_1550_io_x2),
    .io_x3(m_1550_io_x3),
    .io_s(m_1550_io_s),
    .io_cout(m_1550_io_cout)
  );
  Adder m_1551 ( // @[MUL.scala 102:19]
    .io_x1(m_1551_io_x1),
    .io_x2(m_1551_io_x2),
    .io_x3(m_1551_io_x3),
    .io_s(m_1551_io_s),
    .io_cout(m_1551_io_cout)
  );
  Half_Adder m_1552 ( // @[MUL.scala 124:19]
    .io_in_0(m_1552_io_in_0),
    .io_in_1(m_1552_io_in_1),
    .io_out_0(m_1552_io_out_0),
    .io_out_1(m_1552_io_out_1)
  );
  Adder m_1553 ( // @[MUL.scala 102:19]
    .io_x1(m_1553_io_x1),
    .io_x2(m_1553_io_x2),
    .io_x3(m_1553_io_x3),
    .io_s(m_1553_io_s),
    .io_cout(m_1553_io_cout)
  );
  Adder m_1554 ( // @[MUL.scala 102:19]
    .io_x1(m_1554_io_x1),
    .io_x2(m_1554_io_x2),
    .io_x3(m_1554_io_x3),
    .io_s(m_1554_io_s),
    .io_cout(m_1554_io_cout)
  );
  Adder m_1555 ( // @[MUL.scala 102:19]
    .io_x1(m_1555_io_x1),
    .io_x2(m_1555_io_x2),
    .io_x3(m_1555_io_x3),
    .io_s(m_1555_io_s),
    .io_cout(m_1555_io_cout)
  );
  Adder m_1556 ( // @[MUL.scala 102:19]
    .io_x1(m_1556_io_x1),
    .io_x2(m_1556_io_x2),
    .io_x3(m_1556_io_x3),
    .io_s(m_1556_io_s),
    .io_cout(m_1556_io_cout)
  );
  Half_Adder m_1557 ( // @[MUL.scala 124:19]
    .io_in_0(m_1557_io_in_0),
    .io_in_1(m_1557_io_in_1),
    .io_out_0(m_1557_io_out_0),
    .io_out_1(m_1557_io_out_1)
  );
  Adder m_1558 ( // @[MUL.scala 102:19]
    .io_x1(m_1558_io_x1),
    .io_x2(m_1558_io_x2),
    .io_x3(m_1558_io_x3),
    .io_s(m_1558_io_s),
    .io_cout(m_1558_io_cout)
  );
  Adder m_1559 ( // @[MUL.scala 102:19]
    .io_x1(m_1559_io_x1),
    .io_x2(m_1559_io_x2),
    .io_x3(m_1559_io_x3),
    .io_s(m_1559_io_s),
    .io_cout(m_1559_io_cout)
  );
  Adder m_1560 ( // @[MUL.scala 102:19]
    .io_x1(m_1560_io_x1),
    .io_x2(m_1560_io_x2),
    .io_x3(m_1560_io_x3),
    .io_s(m_1560_io_s),
    .io_cout(m_1560_io_cout)
  );
  Adder m_1561 ( // @[MUL.scala 102:19]
    .io_x1(m_1561_io_x1),
    .io_x2(m_1561_io_x2),
    .io_x3(m_1561_io_x3),
    .io_s(m_1561_io_s),
    .io_cout(m_1561_io_cout)
  );
  Half_Adder m_1562 ( // @[MUL.scala 124:19]
    .io_in_0(m_1562_io_in_0),
    .io_in_1(m_1562_io_in_1),
    .io_out_0(m_1562_io_out_0),
    .io_out_1(m_1562_io_out_1)
  );
  Adder m_1563 ( // @[MUL.scala 102:19]
    .io_x1(m_1563_io_x1),
    .io_x2(m_1563_io_x2),
    .io_x3(m_1563_io_x3),
    .io_s(m_1563_io_s),
    .io_cout(m_1563_io_cout)
  );
  Adder m_1564 ( // @[MUL.scala 102:19]
    .io_x1(m_1564_io_x1),
    .io_x2(m_1564_io_x2),
    .io_x3(m_1564_io_x3),
    .io_s(m_1564_io_s),
    .io_cout(m_1564_io_cout)
  );
  Adder m_1565 ( // @[MUL.scala 102:19]
    .io_x1(m_1565_io_x1),
    .io_x2(m_1565_io_x2),
    .io_x3(m_1565_io_x3),
    .io_s(m_1565_io_s),
    .io_cout(m_1565_io_cout)
  );
  Adder m_1566 ( // @[MUL.scala 102:19]
    .io_x1(m_1566_io_x1),
    .io_x2(m_1566_io_x2),
    .io_x3(m_1566_io_x3),
    .io_s(m_1566_io_s),
    .io_cout(m_1566_io_cout)
  );
  Half_Adder m_1567 ( // @[MUL.scala 124:19]
    .io_in_0(m_1567_io_in_0),
    .io_in_1(m_1567_io_in_1),
    .io_out_0(m_1567_io_out_0),
    .io_out_1(m_1567_io_out_1)
  );
  Adder m_1568 ( // @[MUL.scala 102:19]
    .io_x1(m_1568_io_x1),
    .io_x2(m_1568_io_x2),
    .io_x3(m_1568_io_x3),
    .io_s(m_1568_io_s),
    .io_cout(m_1568_io_cout)
  );
  Adder m_1569 ( // @[MUL.scala 102:19]
    .io_x1(m_1569_io_x1),
    .io_x2(m_1569_io_x2),
    .io_x3(m_1569_io_x3),
    .io_s(m_1569_io_s),
    .io_cout(m_1569_io_cout)
  );
  Adder m_1570 ( // @[MUL.scala 102:19]
    .io_x1(m_1570_io_x1),
    .io_x2(m_1570_io_x2),
    .io_x3(m_1570_io_x3),
    .io_s(m_1570_io_s),
    .io_cout(m_1570_io_cout)
  );
  Adder m_1571 ( // @[MUL.scala 102:19]
    .io_x1(m_1571_io_x1),
    .io_x2(m_1571_io_x2),
    .io_x3(m_1571_io_x3),
    .io_s(m_1571_io_s),
    .io_cout(m_1571_io_cout)
  );
  Half_Adder m_1572 ( // @[MUL.scala 124:19]
    .io_in_0(m_1572_io_in_0),
    .io_in_1(m_1572_io_in_1),
    .io_out_0(m_1572_io_out_0),
    .io_out_1(m_1572_io_out_1)
  );
  Adder m_1573 ( // @[MUL.scala 102:19]
    .io_x1(m_1573_io_x1),
    .io_x2(m_1573_io_x2),
    .io_x3(m_1573_io_x3),
    .io_s(m_1573_io_s),
    .io_cout(m_1573_io_cout)
  );
  Adder m_1574 ( // @[MUL.scala 102:19]
    .io_x1(m_1574_io_x1),
    .io_x2(m_1574_io_x2),
    .io_x3(m_1574_io_x3),
    .io_s(m_1574_io_s),
    .io_cout(m_1574_io_cout)
  );
  Adder m_1575 ( // @[MUL.scala 102:19]
    .io_x1(m_1575_io_x1),
    .io_x2(m_1575_io_x2),
    .io_x3(m_1575_io_x3),
    .io_s(m_1575_io_s),
    .io_cout(m_1575_io_cout)
  );
  Adder m_1576 ( // @[MUL.scala 102:19]
    .io_x1(m_1576_io_x1),
    .io_x2(m_1576_io_x2),
    .io_x3(m_1576_io_x3),
    .io_s(m_1576_io_s),
    .io_cout(m_1576_io_cout)
  );
  Adder m_1577 ( // @[MUL.scala 102:19]
    .io_x1(m_1577_io_x1),
    .io_x2(m_1577_io_x2),
    .io_x3(m_1577_io_x3),
    .io_s(m_1577_io_s),
    .io_cout(m_1577_io_cout)
  );
  Adder m_1578 ( // @[MUL.scala 102:19]
    .io_x1(m_1578_io_x1),
    .io_x2(m_1578_io_x2),
    .io_x3(m_1578_io_x3),
    .io_s(m_1578_io_s),
    .io_cout(m_1578_io_cout)
  );
  Adder m_1579 ( // @[MUL.scala 102:19]
    .io_x1(m_1579_io_x1),
    .io_x2(m_1579_io_x2),
    .io_x3(m_1579_io_x3),
    .io_s(m_1579_io_s),
    .io_cout(m_1579_io_cout)
  );
  Adder m_1580 ( // @[MUL.scala 102:19]
    .io_x1(m_1580_io_x1),
    .io_x2(m_1580_io_x2),
    .io_x3(m_1580_io_x3),
    .io_s(m_1580_io_s),
    .io_cout(m_1580_io_cout)
  );
  Adder m_1581 ( // @[MUL.scala 102:19]
    .io_x1(m_1581_io_x1),
    .io_x2(m_1581_io_x2),
    .io_x3(m_1581_io_x3),
    .io_s(m_1581_io_s),
    .io_cout(m_1581_io_cout)
  );
  Adder m_1582 ( // @[MUL.scala 102:19]
    .io_x1(m_1582_io_x1),
    .io_x2(m_1582_io_x2),
    .io_x3(m_1582_io_x3),
    .io_s(m_1582_io_s),
    .io_cout(m_1582_io_cout)
  );
  Adder m_1583 ( // @[MUL.scala 102:19]
    .io_x1(m_1583_io_x1),
    .io_x2(m_1583_io_x2),
    .io_x3(m_1583_io_x3),
    .io_s(m_1583_io_s),
    .io_cout(m_1583_io_cout)
  );
  Adder m_1584 ( // @[MUL.scala 102:19]
    .io_x1(m_1584_io_x1),
    .io_x2(m_1584_io_x2),
    .io_x3(m_1584_io_x3),
    .io_s(m_1584_io_s),
    .io_cout(m_1584_io_cout)
  );
  Adder m_1585 ( // @[MUL.scala 102:19]
    .io_x1(m_1585_io_x1),
    .io_x2(m_1585_io_x2),
    .io_x3(m_1585_io_x3),
    .io_s(m_1585_io_s),
    .io_cout(m_1585_io_cout)
  );
  Adder m_1586 ( // @[MUL.scala 102:19]
    .io_x1(m_1586_io_x1),
    .io_x2(m_1586_io_x2),
    .io_x3(m_1586_io_x3),
    .io_s(m_1586_io_s),
    .io_cout(m_1586_io_cout)
  );
  Adder m_1587 ( // @[MUL.scala 102:19]
    .io_x1(m_1587_io_x1),
    .io_x2(m_1587_io_x2),
    .io_x3(m_1587_io_x3),
    .io_s(m_1587_io_s),
    .io_cout(m_1587_io_cout)
  );
  Adder m_1588 ( // @[MUL.scala 102:19]
    .io_x1(m_1588_io_x1),
    .io_x2(m_1588_io_x2),
    .io_x3(m_1588_io_x3),
    .io_s(m_1588_io_s),
    .io_cout(m_1588_io_cout)
  );
  Adder m_1589 ( // @[MUL.scala 102:19]
    .io_x1(m_1589_io_x1),
    .io_x2(m_1589_io_x2),
    .io_x3(m_1589_io_x3),
    .io_s(m_1589_io_s),
    .io_cout(m_1589_io_cout)
  );
  Adder m_1590 ( // @[MUL.scala 102:19]
    .io_x1(m_1590_io_x1),
    .io_x2(m_1590_io_x2),
    .io_x3(m_1590_io_x3),
    .io_s(m_1590_io_s),
    .io_cout(m_1590_io_cout)
  );
  Adder m_1591 ( // @[MUL.scala 102:19]
    .io_x1(m_1591_io_x1),
    .io_x2(m_1591_io_x2),
    .io_x3(m_1591_io_x3),
    .io_s(m_1591_io_s),
    .io_cout(m_1591_io_cout)
  );
  Adder m_1592 ( // @[MUL.scala 102:19]
    .io_x1(m_1592_io_x1),
    .io_x2(m_1592_io_x2),
    .io_x3(m_1592_io_x3),
    .io_s(m_1592_io_s),
    .io_cout(m_1592_io_cout)
  );
  Adder m_1593 ( // @[MUL.scala 102:19]
    .io_x1(m_1593_io_x1),
    .io_x2(m_1593_io_x2),
    .io_x3(m_1593_io_x3),
    .io_s(m_1593_io_s),
    .io_cout(m_1593_io_cout)
  );
  Adder m_1594 ( // @[MUL.scala 102:19]
    .io_x1(m_1594_io_x1),
    .io_x2(m_1594_io_x2),
    .io_x3(m_1594_io_x3),
    .io_s(m_1594_io_s),
    .io_cout(m_1594_io_cout)
  );
  Adder m_1595 ( // @[MUL.scala 102:19]
    .io_x1(m_1595_io_x1),
    .io_x2(m_1595_io_x2),
    .io_x3(m_1595_io_x3),
    .io_s(m_1595_io_s),
    .io_cout(m_1595_io_cout)
  );
  Adder m_1596 ( // @[MUL.scala 102:19]
    .io_x1(m_1596_io_x1),
    .io_x2(m_1596_io_x2),
    .io_x3(m_1596_io_x3),
    .io_s(m_1596_io_s),
    .io_cout(m_1596_io_cout)
  );
  Adder m_1597 ( // @[MUL.scala 102:19]
    .io_x1(m_1597_io_x1),
    .io_x2(m_1597_io_x2),
    .io_x3(m_1597_io_x3),
    .io_s(m_1597_io_s),
    .io_cout(m_1597_io_cout)
  );
  Adder m_1598 ( // @[MUL.scala 102:19]
    .io_x1(m_1598_io_x1),
    .io_x2(m_1598_io_x2),
    .io_x3(m_1598_io_x3),
    .io_s(m_1598_io_s),
    .io_cout(m_1598_io_cout)
  );
  Adder m_1599 ( // @[MUL.scala 102:19]
    .io_x1(m_1599_io_x1),
    .io_x2(m_1599_io_x2),
    .io_x3(m_1599_io_x3),
    .io_s(m_1599_io_s),
    .io_cout(m_1599_io_cout)
  );
  Adder m_1600 ( // @[MUL.scala 102:19]
    .io_x1(m_1600_io_x1),
    .io_x2(m_1600_io_x2),
    .io_x3(m_1600_io_x3),
    .io_s(m_1600_io_s),
    .io_cout(m_1600_io_cout)
  );
  Adder m_1601 ( // @[MUL.scala 102:19]
    .io_x1(m_1601_io_x1),
    .io_x2(m_1601_io_x2),
    .io_x3(m_1601_io_x3),
    .io_s(m_1601_io_s),
    .io_cout(m_1601_io_cout)
  );
  Adder m_1602 ( // @[MUL.scala 102:19]
    .io_x1(m_1602_io_x1),
    .io_x2(m_1602_io_x2),
    .io_x3(m_1602_io_x3),
    .io_s(m_1602_io_s),
    .io_cout(m_1602_io_cout)
  );
  Adder m_1603 ( // @[MUL.scala 102:19]
    .io_x1(m_1603_io_x1),
    .io_x2(m_1603_io_x2),
    .io_x3(m_1603_io_x3),
    .io_s(m_1603_io_s),
    .io_cout(m_1603_io_cout)
  );
  Half_Adder m_1604 ( // @[MUL.scala 124:19]
    .io_in_0(m_1604_io_in_0),
    .io_in_1(m_1604_io_in_1),
    .io_out_0(m_1604_io_out_0),
    .io_out_1(m_1604_io_out_1)
  );
  Adder m_1605 ( // @[MUL.scala 102:19]
    .io_x1(m_1605_io_x1),
    .io_x2(m_1605_io_x2),
    .io_x3(m_1605_io_x3),
    .io_s(m_1605_io_s),
    .io_cout(m_1605_io_cout)
  );
  Adder m_1606 ( // @[MUL.scala 102:19]
    .io_x1(m_1606_io_x1),
    .io_x2(m_1606_io_x2),
    .io_x3(m_1606_io_x3),
    .io_s(m_1606_io_s),
    .io_cout(m_1606_io_cout)
  );
  Adder m_1607 ( // @[MUL.scala 102:19]
    .io_x1(m_1607_io_x1),
    .io_x2(m_1607_io_x2),
    .io_x3(m_1607_io_x3),
    .io_s(m_1607_io_s),
    .io_cout(m_1607_io_cout)
  );
  Half_Adder m_1608 ( // @[MUL.scala 124:19]
    .io_in_0(m_1608_io_in_0),
    .io_in_1(m_1608_io_in_1),
    .io_out_0(m_1608_io_out_0),
    .io_out_1(m_1608_io_out_1)
  );
  Adder m_1609 ( // @[MUL.scala 102:19]
    .io_x1(m_1609_io_x1),
    .io_x2(m_1609_io_x2),
    .io_x3(m_1609_io_x3),
    .io_s(m_1609_io_s),
    .io_cout(m_1609_io_cout)
  );
  Adder m_1610 ( // @[MUL.scala 102:19]
    .io_x1(m_1610_io_x1),
    .io_x2(m_1610_io_x2),
    .io_x3(m_1610_io_x3),
    .io_s(m_1610_io_s),
    .io_cout(m_1610_io_cout)
  );
  Adder m_1611 ( // @[MUL.scala 102:19]
    .io_x1(m_1611_io_x1),
    .io_x2(m_1611_io_x2),
    .io_x3(m_1611_io_x3),
    .io_s(m_1611_io_s),
    .io_cout(m_1611_io_cout)
  );
  Half_Adder m_1612 ( // @[MUL.scala 124:19]
    .io_in_0(m_1612_io_in_0),
    .io_in_1(m_1612_io_in_1),
    .io_out_0(m_1612_io_out_0),
    .io_out_1(m_1612_io_out_1)
  );
  Adder m_1613 ( // @[MUL.scala 102:19]
    .io_x1(m_1613_io_x1),
    .io_x2(m_1613_io_x2),
    .io_x3(m_1613_io_x3),
    .io_s(m_1613_io_s),
    .io_cout(m_1613_io_cout)
  );
  Adder m_1614 ( // @[MUL.scala 102:19]
    .io_x1(m_1614_io_x1),
    .io_x2(m_1614_io_x2),
    .io_x3(m_1614_io_x3),
    .io_s(m_1614_io_s),
    .io_cout(m_1614_io_cout)
  );
  Adder m_1615 ( // @[MUL.scala 102:19]
    .io_x1(m_1615_io_x1),
    .io_x2(m_1615_io_x2),
    .io_x3(m_1615_io_x3),
    .io_s(m_1615_io_s),
    .io_cout(m_1615_io_cout)
  );
  Half_Adder m_1616 ( // @[MUL.scala 124:19]
    .io_in_0(m_1616_io_in_0),
    .io_in_1(m_1616_io_in_1),
    .io_out_0(m_1616_io_out_0),
    .io_out_1(m_1616_io_out_1)
  );
  Adder m_1617 ( // @[MUL.scala 102:19]
    .io_x1(m_1617_io_x1),
    .io_x2(m_1617_io_x2),
    .io_x3(m_1617_io_x3),
    .io_s(m_1617_io_s),
    .io_cout(m_1617_io_cout)
  );
  Adder m_1618 ( // @[MUL.scala 102:19]
    .io_x1(m_1618_io_x1),
    .io_x2(m_1618_io_x2),
    .io_x3(m_1618_io_x3),
    .io_s(m_1618_io_s),
    .io_cout(m_1618_io_cout)
  );
  Adder m_1619 ( // @[MUL.scala 102:19]
    .io_x1(m_1619_io_x1),
    .io_x2(m_1619_io_x2),
    .io_x3(m_1619_io_x3),
    .io_s(m_1619_io_s),
    .io_cout(m_1619_io_cout)
  );
  Adder m_1620 ( // @[MUL.scala 102:19]
    .io_x1(m_1620_io_x1),
    .io_x2(m_1620_io_x2),
    .io_x3(m_1620_io_x3),
    .io_s(m_1620_io_s),
    .io_cout(m_1620_io_cout)
  );
  Adder m_1621 ( // @[MUL.scala 102:19]
    .io_x1(m_1621_io_x1),
    .io_x2(m_1621_io_x2),
    .io_x3(m_1621_io_x3),
    .io_s(m_1621_io_s),
    .io_cout(m_1621_io_cout)
  );
  Adder m_1622 ( // @[MUL.scala 102:19]
    .io_x1(m_1622_io_x1),
    .io_x2(m_1622_io_x2),
    .io_x3(m_1622_io_x3),
    .io_s(m_1622_io_s),
    .io_cout(m_1622_io_cout)
  );
  Adder m_1623 ( // @[MUL.scala 102:19]
    .io_x1(m_1623_io_x1),
    .io_x2(m_1623_io_x2),
    .io_x3(m_1623_io_x3),
    .io_s(m_1623_io_s),
    .io_cout(m_1623_io_cout)
  );
  Adder m_1624 ( // @[MUL.scala 102:19]
    .io_x1(m_1624_io_x1),
    .io_x2(m_1624_io_x2),
    .io_x3(m_1624_io_x3),
    .io_s(m_1624_io_s),
    .io_cout(m_1624_io_cout)
  );
  Adder m_1625 ( // @[MUL.scala 102:19]
    .io_x1(m_1625_io_x1),
    .io_x2(m_1625_io_x2),
    .io_x3(m_1625_io_x3),
    .io_s(m_1625_io_s),
    .io_cout(m_1625_io_cout)
  );
  Adder m_1626 ( // @[MUL.scala 102:19]
    .io_x1(m_1626_io_x1),
    .io_x2(m_1626_io_x2),
    .io_x3(m_1626_io_x3),
    .io_s(m_1626_io_s),
    .io_cout(m_1626_io_cout)
  );
  Adder m_1627 ( // @[MUL.scala 102:19]
    .io_x1(m_1627_io_x1),
    .io_x2(m_1627_io_x2),
    .io_x3(m_1627_io_x3),
    .io_s(m_1627_io_s),
    .io_cout(m_1627_io_cout)
  );
  Adder m_1628 ( // @[MUL.scala 102:19]
    .io_x1(m_1628_io_x1),
    .io_x2(m_1628_io_x2),
    .io_x3(m_1628_io_x3),
    .io_s(m_1628_io_s),
    .io_cout(m_1628_io_cout)
  );
  Adder m_1629 ( // @[MUL.scala 102:19]
    .io_x1(m_1629_io_x1),
    .io_x2(m_1629_io_x2),
    .io_x3(m_1629_io_x3),
    .io_s(m_1629_io_s),
    .io_cout(m_1629_io_cout)
  );
  Adder m_1630 ( // @[MUL.scala 102:19]
    .io_x1(m_1630_io_x1),
    .io_x2(m_1630_io_x2),
    .io_x3(m_1630_io_x3),
    .io_s(m_1630_io_s),
    .io_cout(m_1630_io_cout)
  );
  Adder m_1631 ( // @[MUL.scala 102:19]
    .io_x1(m_1631_io_x1),
    .io_x2(m_1631_io_x2),
    .io_x3(m_1631_io_x3),
    .io_s(m_1631_io_s),
    .io_cout(m_1631_io_cout)
  );
  Adder m_1632 ( // @[MUL.scala 102:19]
    .io_x1(m_1632_io_x1),
    .io_x2(m_1632_io_x2),
    .io_x3(m_1632_io_x3),
    .io_s(m_1632_io_s),
    .io_cout(m_1632_io_cout)
  );
  Adder m_1633 ( // @[MUL.scala 102:19]
    .io_x1(m_1633_io_x1),
    .io_x2(m_1633_io_x2),
    .io_x3(m_1633_io_x3),
    .io_s(m_1633_io_s),
    .io_cout(m_1633_io_cout)
  );
  Adder m_1634 ( // @[MUL.scala 102:19]
    .io_x1(m_1634_io_x1),
    .io_x2(m_1634_io_x2),
    .io_x3(m_1634_io_x3),
    .io_s(m_1634_io_s),
    .io_cout(m_1634_io_cout)
  );
  Adder m_1635 ( // @[MUL.scala 102:19]
    .io_x1(m_1635_io_x1),
    .io_x2(m_1635_io_x2),
    .io_x3(m_1635_io_x3),
    .io_s(m_1635_io_s),
    .io_cout(m_1635_io_cout)
  );
  Adder m_1636 ( // @[MUL.scala 102:19]
    .io_x1(m_1636_io_x1),
    .io_x2(m_1636_io_x2),
    .io_x3(m_1636_io_x3),
    .io_s(m_1636_io_s),
    .io_cout(m_1636_io_cout)
  );
  Adder m_1637 ( // @[MUL.scala 102:19]
    .io_x1(m_1637_io_x1),
    .io_x2(m_1637_io_x2),
    .io_x3(m_1637_io_x3),
    .io_s(m_1637_io_s),
    .io_cout(m_1637_io_cout)
  );
  Adder m_1638 ( // @[MUL.scala 102:19]
    .io_x1(m_1638_io_x1),
    .io_x2(m_1638_io_x2),
    .io_x3(m_1638_io_x3),
    .io_s(m_1638_io_s),
    .io_cout(m_1638_io_cout)
  );
  Adder m_1639 ( // @[MUL.scala 102:19]
    .io_x1(m_1639_io_x1),
    .io_x2(m_1639_io_x2),
    .io_x3(m_1639_io_x3),
    .io_s(m_1639_io_s),
    .io_cout(m_1639_io_cout)
  );
  Half_Adder m_1640 ( // @[MUL.scala 124:19]
    .io_in_0(m_1640_io_in_0),
    .io_in_1(m_1640_io_in_1),
    .io_out_0(m_1640_io_out_0),
    .io_out_1(m_1640_io_out_1)
  );
  Adder m_1641 ( // @[MUL.scala 102:19]
    .io_x1(m_1641_io_x1),
    .io_x2(m_1641_io_x2),
    .io_x3(m_1641_io_x3),
    .io_s(m_1641_io_s),
    .io_cout(m_1641_io_cout)
  );
  Adder m_1642 ( // @[MUL.scala 102:19]
    .io_x1(m_1642_io_x1),
    .io_x2(m_1642_io_x2),
    .io_x3(m_1642_io_x3),
    .io_s(m_1642_io_s),
    .io_cout(m_1642_io_cout)
  );
  Half_Adder m_1643 ( // @[MUL.scala 124:19]
    .io_in_0(m_1643_io_in_0),
    .io_in_1(m_1643_io_in_1),
    .io_out_0(m_1643_io_out_0),
    .io_out_1(m_1643_io_out_1)
  );
  Adder m_1644 ( // @[MUL.scala 102:19]
    .io_x1(m_1644_io_x1),
    .io_x2(m_1644_io_x2),
    .io_x3(m_1644_io_x3),
    .io_s(m_1644_io_s),
    .io_cout(m_1644_io_cout)
  );
  Adder m_1645 ( // @[MUL.scala 102:19]
    .io_x1(m_1645_io_x1),
    .io_x2(m_1645_io_x2),
    .io_x3(m_1645_io_x3),
    .io_s(m_1645_io_s),
    .io_cout(m_1645_io_cout)
  );
  Half_Adder m_1646 ( // @[MUL.scala 124:19]
    .io_in_0(m_1646_io_in_0),
    .io_in_1(m_1646_io_in_1),
    .io_out_0(m_1646_io_out_0),
    .io_out_1(m_1646_io_out_1)
  );
  Adder m_1647 ( // @[MUL.scala 102:19]
    .io_x1(m_1647_io_x1),
    .io_x2(m_1647_io_x2),
    .io_x3(m_1647_io_x3),
    .io_s(m_1647_io_s),
    .io_cout(m_1647_io_cout)
  );
  Adder m_1648 ( // @[MUL.scala 102:19]
    .io_x1(m_1648_io_x1),
    .io_x2(m_1648_io_x2),
    .io_x3(m_1648_io_x3),
    .io_s(m_1648_io_s),
    .io_cout(m_1648_io_cout)
  );
  Half_Adder m_1649 ( // @[MUL.scala 124:19]
    .io_in_0(m_1649_io_in_0),
    .io_in_1(m_1649_io_in_1),
    .io_out_0(m_1649_io_out_0),
    .io_out_1(m_1649_io_out_1)
  );
  Adder m_1650 ( // @[MUL.scala 102:19]
    .io_x1(m_1650_io_x1),
    .io_x2(m_1650_io_x2),
    .io_x3(m_1650_io_x3),
    .io_s(m_1650_io_s),
    .io_cout(m_1650_io_cout)
  );
  Adder m_1651 ( // @[MUL.scala 102:19]
    .io_x1(m_1651_io_x1),
    .io_x2(m_1651_io_x2),
    .io_x3(m_1651_io_x3),
    .io_s(m_1651_io_s),
    .io_cout(m_1651_io_cout)
  );
  Half_Adder m_1652 ( // @[MUL.scala 124:19]
    .io_in_0(m_1652_io_in_0),
    .io_in_1(m_1652_io_in_1),
    .io_out_0(m_1652_io_out_0),
    .io_out_1(m_1652_io_out_1)
  );
  Adder m_1653 ( // @[MUL.scala 102:19]
    .io_x1(m_1653_io_x1),
    .io_x2(m_1653_io_x2),
    .io_x3(m_1653_io_x3),
    .io_s(m_1653_io_s),
    .io_cout(m_1653_io_cout)
  );
  Adder m_1654 ( // @[MUL.scala 102:19]
    .io_x1(m_1654_io_x1),
    .io_x2(m_1654_io_x2),
    .io_x3(m_1654_io_x3),
    .io_s(m_1654_io_s),
    .io_cout(m_1654_io_cout)
  );
  Half_Adder m_1655 ( // @[MUL.scala 124:19]
    .io_in_0(m_1655_io_in_0),
    .io_in_1(m_1655_io_in_1),
    .io_out_0(m_1655_io_out_0),
    .io_out_1(m_1655_io_out_1)
  );
  Adder m_1656 ( // @[MUL.scala 102:19]
    .io_x1(m_1656_io_x1),
    .io_x2(m_1656_io_x2),
    .io_x3(m_1656_io_x3),
    .io_s(m_1656_io_s),
    .io_cout(m_1656_io_cout)
  );
  Adder m_1657 ( // @[MUL.scala 102:19]
    .io_x1(m_1657_io_x1),
    .io_x2(m_1657_io_x2),
    .io_x3(m_1657_io_x3),
    .io_s(m_1657_io_s),
    .io_cout(m_1657_io_cout)
  );
  Half_Adder m_1658 ( // @[MUL.scala 124:19]
    .io_in_0(m_1658_io_in_0),
    .io_in_1(m_1658_io_in_1),
    .io_out_0(m_1658_io_out_0),
    .io_out_1(m_1658_io_out_1)
  );
  Adder m_1659 ( // @[MUL.scala 102:19]
    .io_x1(m_1659_io_x1),
    .io_x2(m_1659_io_x2),
    .io_x3(m_1659_io_x3),
    .io_s(m_1659_io_s),
    .io_cout(m_1659_io_cout)
  );
  Adder m_1660 ( // @[MUL.scala 102:19]
    .io_x1(m_1660_io_x1),
    .io_x2(m_1660_io_x2),
    .io_x3(m_1660_io_x3),
    .io_s(m_1660_io_s),
    .io_cout(m_1660_io_cout)
  );
  Adder m_1661 ( // @[MUL.scala 102:19]
    .io_x1(m_1661_io_x1),
    .io_x2(m_1661_io_x2),
    .io_x3(m_1661_io_x3),
    .io_s(m_1661_io_s),
    .io_cout(m_1661_io_cout)
  );
  Adder m_1662 ( // @[MUL.scala 102:19]
    .io_x1(m_1662_io_x1),
    .io_x2(m_1662_io_x2),
    .io_x3(m_1662_io_x3),
    .io_s(m_1662_io_s),
    .io_cout(m_1662_io_cout)
  );
  Adder m_1663 ( // @[MUL.scala 102:19]
    .io_x1(m_1663_io_x1),
    .io_x2(m_1663_io_x2),
    .io_x3(m_1663_io_x3),
    .io_s(m_1663_io_s),
    .io_cout(m_1663_io_cout)
  );
  Adder m_1664 ( // @[MUL.scala 102:19]
    .io_x1(m_1664_io_x1),
    .io_x2(m_1664_io_x2),
    .io_x3(m_1664_io_x3),
    .io_s(m_1664_io_s),
    .io_cout(m_1664_io_cout)
  );
  Adder m_1665 ( // @[MUL.scala 102:19]
    .io_x1(m_1665_io_x1),
    .io_x2(m_1665_io_x2),
    .io_x3(m_1665_io_x3),
    .io_s(m_1665_io_s),
    .io_cout(m_1665_io_cout)
  );
  Adder m_1666 ( // @[MUL.scala 102:19]
    .io_x1(m_1666_io_x1),
    .io_x2(m_1666_io_x2),
    .io_x3(m_1666_io_x3),
    .io_s(m_1666_io_s),
    .io_cout(m_1666_io_cout)
  );
  Adder m_1667 ( // @[MUL.scala 102:19]
    .io_x1(m_1667_io_x1),
    .io_x2(m_1667_io_x2),
    .io_x3(m_1667_io_x3),
    .io_s(m_1667_io_s),
    .io_cout(m_1667_io_cout)
  );
  Adder m_1668 ( // @[MUL.scala 102:19]
    .io_x1(m_1668_io_x1),
    .io_x2(m_1668_io_x2),
    .io_x3(m_1668_io_x3),
    .io_s(m_1668_io_s),
    .io_cout(m_1668_io_cout)
  );
  Adder m_1669 ( // @[MUL.scala 102:19]
    .io_x1(m_1669_io_x1),
    .io_x2(m_1669_io_x2),
    .io_x3(m_1669_io_x3),
    .io_s(m_1669_io_s),
    .io_cout(m_1669_io_cout)
  );
  Adder m_1670 ( // @[MUL.scala 102:19]
    .io_x1(m_1670_io_x1),
    .io_x2(m_1670_io_x2),
    .io_x3(m_1670_io_x3),
    .io_s(m_1670_io_s),
    .io_cout(m_1670_io_cout)
  );
  Adder m_1671 ( // @[MUL.scala 102:19]
    .io_x1(m_1671_io_x1),
    .io_x2(m_1671_io_x2),
    .io_x3(m_1671_io_x3),
    .io_s(m_1671_io_s),
    .io_cout(m_1671_io_cout)
  );
  Adder m_1672 ( // @[MUL.scala 102:19]
    .io_x1(m_1672_io_x1),
    .io_x2(m_1672_io_x2),
    .io_x3(m_1672_io_x3),
    .io_s(m_1672_io_s),
    .io_cout(m_1672_io_cout)
  );
  Adder m_1673 ( // @[MUL.scala 102:19]
    .io_x1(m_1673_io_x1),
    .io_x2(m_1673_io_x2),
    .io_x3(m_1673_io_x3),
    .io_s(m_1673_io_s),
    .io_cout(m_1673_io_cout)
  );
  Adder m_1674 ( // @[MUL.scala 102:19]
    .io_x1(m_1674_io_x1),
    .io_x2(m_1674_io_x2),
    .io_x3(m_1674_io_x3),
    .io_s(m_1674_io_s),
    .io_cout(m_1674_io_cout)
  );
  Adder m_1675 ( // @[MUL.scala 102:19]
    .io_x1(m_1675_io_x1),
    .io_x2(m_1675_io_x2),
    .io_x3(m_1675_io_x3),
    .io_s(m_1675_io_s),
    .io_cout(m_1675_io_cout)
  );
  Adder m_1676 ( // @[MUL.scala 102:19]
    .io_x1(m_1676_io_x1),
    .io_x2(m_1676_io_x2),
    .io_x3(m_1676_io_x3),
    .io_s(m_1676_io_s),
    .io_cout(m_1676_io_cout)
  );
  Adder m_1677 ( // @[MUL.scala 102:19]
    .io_x1(m_1677_io_x1),
    .io_x2(m_1677_io_x2),
    .io_x3(m_1677_io_x3),
    .io_s(m_1677_io_s),
    .io_cout(m_1677_io_cout)
  );
  Adder m_1678 ( // @[MUL.scala 102:19]
    .io_x1(m_1678_io_x1),
    .io_x2(m_1678_io_x2),
    .io_x3(m_1678_io_x3),
    .io_s(m_1678_io_s),
    .io_cout(m_1678_io_cout)
  );
  Adder m_1679 ( // @[MUL.scala 102:19]
    .io_x1(m_1679_io_x1),
    .io_x2(m_1679_io_x2),
    .io_x3(m_1679_io_x3),
    .io_s(m_1679_io_s),
    .io_cout(m_1679_io_cout)
  );
  Adder m_1680 ( // @[MUL.scala 102:19]
    .io_x1(m_1680_io_x1),
    .io_x2(m_1680_io_x2),
    .io_x3(m_1680_io_x3),
    .io_s(m_1680_io_s),
    .io_cout(m_1680_io_cout)
  );
  Adder m_1681 ( // @[MUL.scala 102:19]
    .io_x1(m_1681_io_x1),
    .io_x2(m_1681_io_x2),
    .io_x3(m_1681_io_x3),
    .io_s(m_1681_io_s),
    .io_cout(m_1681_io_cout)
  );
  Adder m_1682 ( // @[MUL.scala 102:19]
    .io_x1(m_1682_io_x1),
    .io_x2(m_1682_io_x2),
    .io_x3(m_1682_io_x3),
    .io_s(m_1682_io_s),
    .io_cout(m_1682_io_cout)
  );
  Adder m_1683 ( // @[MUL.scala 102:19]
    .io_x1(m_1683_io_x1),
    .io_x2(m_1683_io_x2),
    .io_x3(m_1683_io_x3),
    .io_s(m_1683_io_s),
    .io_cout(m_1683_io_cout)
  );
  Adder m_1684 ( // @[MUL.scala 102:19]
    .io_x1(m_1684_io_x1),
    .io_x2(m_1684_io_x2),
    .io_x3(m_1684_io_x3),
    .io_s(m_1684_io_s),
    .io_cout(m_1684_io_cout)
  );
  Adder m_1685 ( // @[MUL.scala 102:19]
    .io_x1(m_1685_io_x1),
    .io_x2(m_1685_io_x2),
    .io_x3(m_1685_io_x3),
    .io_s(m_1685_io_s),
    .io_cout(m_1685_io_cout)
  );
  Adder m_1686 ( // @[MUL.scala 102:19]
    .io_x1(m_1686_io_x1),
    .io_x2(m_1686_io_x2),
    .io_x3(m_1686_io_x3),
    .io_s(m_1686_io_s),
    .io_cout(m_1686_io_cout)
  );
  Adder m_1687 ( // @[MUL.scala 102:19]
    .io_x1(m_1687_io_x1),
    .io_x2(m_1687_io_x2),
    .io_x3(m_1687_io_x3),
    .io_s(m_1687_io_s),
    .io_cout(m_1687_io_cout)
  );
  Adder m_1688 ( // @[MUL.scala 102:19]
    .io_x1(m_1688_io_x1),
    .io_x2(m_1688_io_x2),
    .io_x3(m_1688_io_x3),
    .io_s(m_1688_io_s),
    .io_cout(m_1688_io_cout)
  );
  Adder m_1689 ( // @[MUL.scala 102:19]
    .io_x1(m_1689_io_x1),
    .io_x2(m_1689_io_x2),
    .io_x3(m_1689_io_x3),
    .io_s(m_1689_io_s),
    .io_cout(m_1689_io_cout)
  );
  Adder m_1690 ( // @[MUL.scala 102:19]
    .io_x1(m_1690_io_x1),
    .io_x2(m_1690_io_x2),
    .io_x3(m_1690_io_x3),
    .io_s(m_1690_io_s),
    .io_cout(m_1690_io_cout)
  );
  Adder m_1691 ( // @[MUL.scala 102:19]
    .io_x1(m_1691_io_x1),
    .io_x2(m_1691_io_x2),
    .io_x3(m_1691_io_x3),
    .io_s(m_1691_io_s),
    .io_cout(m_1691_io_cout)
  );
  Half_Adder m_1692 ( // @[MUL.scala 124:19]
    .io_in_0(m_1692_io_in_0),
    .io_in_1(m_1692_io_in_1),
    .io_out_0(m_1692_io_out_0),
    .io_out_1(m_1692_io_out_1)
  );
  Half_Adder m_1693 ( // @[MUL.scala 124:19]
    .io_in_0(m_1693_io_in_0),
    .io_in_1(m_1693_io_in_1),
    .io_out_0(m_1693_io_out_0),
    .io_out_1(m_1693_io_out_1)
  );
  Half_Adder m_1694 ( // @[MUL.scala 124:19]
    .io_in_0(m_1694_io_in_0),
    .io_in_1(m_1694_io_in_1),
    .io_out_0(m_1694_io_out_0),
    .io_out_1(m_1694_io_out_1)
  );
  Half_Adder m_1695 ( // @[MUL.scala 124:19]
    .io_in_0(m_1695_io_in_0),
    .io_in_1(m_1695_io_in_1),
    .io_out_0(m_1695_io_out_0),
    .io_out_1(m_1695_io_out_1)
  );
  Half_Adder m_1696 ( // @[MUL.scala 124:19]
    .io_in_0(m_1696_io_in_0),
    .io_in_1(m_1696_io_in_1),
    .io_out_0(m_1696_io_out_0),
    .io_out_1(m_1696_io_out_1)
  );
  Half_Adder m_1697 ( // @[MUL.scala 124:19]
    .io_in_0(m_1697_io_in_0),
    .io_in_1(m_1697_io_in_1),
    .io_out_0(m_1697_io_out_0),
    .io_out_1(m_1697_io_out_1)
  );
  Half_Adder m_1698 ( // @[MUL.scala 124:19]
    .io_in_0(m_1698_io_in_0),
    .io_in_1(m_1698_io_in_1),
    .io_out_0(m_1698_io_out_0),
    .io_out_1(m_1698_io_out_1)
  );
  Half_Adder m_1699 ( // @[MUL.scala 124:19]
    .io_in_0(m_1699_io_in_0),
    .io_in_1(m_1699_io_in_1),
    .io_out_0(m_1699_io_out_0),
    .io_out_1(m_1699_io_out_1)
  );
  Half_Adder m_1700 ( // @[MUL.scala 124:19]
    .io_in_0(m_1700_io_in_0),
    .io_in_1(m_1700_io_in_1),
    .io_out_0(m_1700_io_out_0),
    .io_out_1(m_1700_io_out_1)
  );
  Half_Adder m_1701 ( // @[MUL.scala 124:19]
    .io_in_0(m_1701_io_in_0),
    .io_in_1(m_1701_io_in_1),
    .io_out_0(m_1701_io_out_0),
    .io_out_1(m_1701_io_out_1)
  );
  Half_Adder m_1702 ( // @[MUL.scala 124:19]
    .io_in_0(m_1702_io_in_0),
    .io_in_1(m_1702_io_in_1),
    .io_out_0(m_1702_io_out_0),
    .io_out_1(m_1702_io_out_1)
  );
  Half_Adder m_1703 ( // @[MUL.scala 124:19]
    .io_in_0(m_1703_io_in_0),
    .io_in_1(m_1703_io_in_1),
    .io_out_0(m_1703_io_out_0),
    .io_out_1(m_1703_io_out_1)
  );
  Half_Adder m_1704 ( // @[MUL.scala 124:19]
    .io_in_0(m_1704_io_in_0),
    .io_in_1(m_1704_io_in_1),
    .io_out_0(m_1704_io_out_0),
    .io_out_1(m_1704_io_out_1)
  );
  Half_Adder m_1705 ( // @[MUL.scala 124:19]
    .io_in_0(m_1705_io_in_0),
    .io_in_1(m_1705_io_in_1),
    .io_out_0(m_1705_io_out_0),
    .io_out_1(m_1705_io_out_1)
  );
  Adder m_1706 ( // @[MUL.scala 102:19]
    .io_x1(m_1706_io_x1),
    .io_x2(m_1706_io_x2),
    .io_x3(m_1706_io_x3),
    .io_s(m_1706_io_s),
    .io_cout(m_1706_io_cout)
  );
  Adder m_1707 ( // @[MUL.scala 102:19]
    .io_x1(m_1707_io_x1),
    .io_x2(m_1707_io_x2),
    .io_x3(m_1707_io_x3),
    .io_s(m_1707_io_s),
    .io_cout(m_1707_io_cout)
  );
  Adder m_1708 ( // @[MUL.scala 102:19]
    .io_x1(m_1708_io_x1),
    .io_x2(m_1708_io_x2),
    .io_x3(m_1708_io_x3),
    .io_s(m_1708_io_s),
    .io_cout(m_1708_io_cout)
  );
  Adder m_1709 ( // @[MUL.scala 102:19]
    .io_x1(m_1709_io_x1),
    .io_x2(m_1709_io_x2),
    .io_x3(m_1709_io_x3),
    .io_s(m_1709_io_s),
    .io_cout(m_1709_io_cout)
  );
  Adder m_1710 ( // @[MUL.scala 102:19]
    .io_x1(m_1710_io_x1),
    .io_x2(m_1710_io_x2),
    .io_x3(m_1710_io_x3),
    .io_s(m_1710_io_s),
    .io_cout(m_1710_io_cout)
  );
  Adder m_1711 ( // @[MUL.scala 102:19]
    .io_x1(m_1711_io_x1),
    .io_x2(m_1711_io_x2),
    .io_x3(m_1711_io_x3),
    .io_s(m_1711_io_s),
    .io_cout(m_1711_io_cout)
  );
  Adder m_1712 ( // @[MUL.scala 102:19]
    .io_x1(m_1712_io_x1),
    .io_x2(m_1712_io_x2),
    .io_x3(m_1712_io_x3),
    .io_s(m_1712_io_s),
    .io_cout(m_1712_io_cout)
  );
  Adder m_1713 ( // @[MUL.scala 102:19]
    .io_x1(m_1713_io_x1),
    .io_x2(m_1713_io_x2),
    .io_x3(m_1713_io_x3),
    .io_s(m_1713_io_s),
    .io_cout(m_1713_io_cout)
  );
  Adder m_1714 ( // @[MUL.scala 102:19]
    .io_x1(m_1714_io_x1),
    .io_x2(m_1714_io_x2),
    .io_x3(m_1714_io_x3),
    .io_s(m_1714_io_s),
    .io_cout(m_1714_io_cout)
  );
  Adder m_1715 ( // @[MUL.scala 102:19]
    .io_x1(m_1715_io_x1),
    .io_x2(m_1715_io_x2),
    .io_x3(m_1715_io_x3),
    .io_s(m_1715_io_s),
    .io_cout(m_1715_io_cout)
  );
  Adder m_1716 ( // @[MUL.scala 102:19]
    .io_x1(m_1716_io_x1),
    .io_x2(m_1716_io_x2),
    .io_x3(m_1716_io_x3),
    .io_s(m_1716_io_s),
    .io_cout(m_1716_io_cout)
  );
  Adder m_1717 ( // @[MUL.scala 102:19]
    .io_x1(m_1717_io_x1),
    .io_x2(m_1717_io_x2),
    .io_x3(m_1717_io_x3),
    .io_s(m_1717_io_s),
    .io_cout(m_1717_io_cout)
  );
  Adder m_1718 ( // @[MUL.scala 102:19]
    .io_x1(m_1718_io_x1),
    .io_x2(m_1718_io_x2),
    .io_x3(m_1718_io_x3),
    .io_s(m_1718_io_s),
    .io_cout(m_1718_io_cout)
  );
  Adder m_1719 ( // @[MUL.scala 102:19]
    .io_x1(m_1719_io_x1),
    .io_x2(m_1719_io_x2),
    .io_x3(m_1719_io_x3),
    .io_s(m_1719_io_s),
    .io_cout(m_1719_io_cout)
  );
  Adder m_1720 ( // @[MUL.scala 102:19]
    .io_x1(m_1720_io_x1),
    .io_x2(m_1720_io_x2),
    .io_x3(m_1720_io_x3),
    .io_s(m_1720_io_s),
    .io_cout(m_1720_io_cout)
  );
  Half_Adder m_1721 ( // @[MUL.scala 124:19]
    .io_in_0(m_1721_io_in_0),
    .io_in_1(m_1721_io_in_1),
    .io_out_0(m_1721_io_out_0),
    .io_out_1(m_1721_io_out_1)
  );
  Adder m_1722 ( // @[MUL.scala 102:19]
    .io_x1(m_1722_io_x1),
    .io_x2(m_1722_io_x2),
    .io_x3(m_1722_io_x3),
    .io_s(m_1722_io_s),
    .io_cout(m_1722_io_cout)
  );
  Half_Adder m_1723 ( // @[MUL.scala 124:19]
    .io_in_0(m_1723_io_in_0),
    .io_in_1(m_1723_io_in_1),
    .io_out_0(m_1723_io_out_0),
    .io_out_1(m_1723_io_out_1)
  );
  Adder m_1724 ( // @[MUL.scala 102:19]
    .io_x1(m_1724_io_x1),
    .io_x2(m_1724_io_x2),
    .io_x3(m_1724_io_x3),
    .io_s(m_1724_io_s),
    .io_cout(m_1724_io_cout)
  );
  Half_Adder m_1725 ( // @[MUL.scala 124:19]
    .io_in_0(m_1725_io_in_0),
    .io_in_1(m_1725_io_in_1),
    .io_out_0(m_1725_io_out_0),
    .io_out_1(m_1725_io_out_1)
  );
  Adder m_1726 ( // @[MUL.scala 102:19]
    .io_x1(m_1726_io_x1),
    .io_x2(m_1726_io_x2),
    .io_x3(m_1726_io_x3),
    .io_s(m_1726_io_s),
    .io_cout(m_1726_io_cout)
  );
  Half_Adder m_1727 ( // @[MUL.scala 124:19]
    .io_in_0(m_1727_io_in_0),
    .io_in_1(m_1727_io_in_1),
    .io_out_0(m_1727_io_out_0),
    .io_out_1(m_1727_io_out_1)
  );
  Adder m_1728 ( // @[MUL.scala 102:19]
    .io_x1(m_1728_io_x1),
    .io_x2(m_1728_io_x2),
    .io_x3(m_1728_io_x3),
    .io_s(m_1728_io_s),
    .io_cout(m_1728_io_cout)
  );
  Half_Adder m_1729 ( // @[MUL.scala 124:19]
    .io_in_0(m_1729_io_in_0),
    .io_in_1(m_1729_io_in_1),
    .io_out_0(m_1729_io_out_0),
    .io_out_1(m_1729_io_out_1)
  );
  Adder m_1730 ( // @[MUL.scala 102:19]
    .io_x1(m_1730_io_x1),
    .io_x2(m_1730_io_x2),
    .io_x3(m_1730_io_x3),
    .io_s(m_1730_io_s),
    .io_cout(m_1730_io_cout)
  );
  Adder m_1731 ( // @[MUL.scala 102:19]
    .io_x1(m_1731_io_x1),
    .io_x2(m_1731_io_x2),
    .io_x3(m_1731_io_x3),
    .io_s(m_1731_io_s),
    .io_cout(m_1731_io_cout)
  );
  Adder m_1732 ( // @[MUL.scala 102:19]
    .io_x1(m_1732_io_x1),
    .io_x2(m_1732_io_x2),
    .io_x3(m_1732_io_x3),
    .io_s(m_1732_io_s),
    .io_cout(m_1732_io_cout)
  );
  Adder m_1733 ( // @[MUL.scala 102:19]
    .io_x1(m_1733_io_x1),
    .io_x2(m_1733_io_x2),
    .io_x3(m_1733_io_x3),
    .io_s(m_1733_io_s),
    .io_cout(m_1733_io_cout)
  );
  Adder m_1734 ( // @[MUL.scala 102:19]
    .io_x1(m_1734_io_x1),
    .io_x2(m_1734_io_x2),
    .io_x3(m_1734_io_x3),
    .io_s(m_1734_io_s),
    .io_cout(m_1734_io_cout)
  );
  Adder m_1735 ( // @[MUL.scala 102:19]
    .io_x1(m_1735_io_x1),
    .io_x2(m_1735_io_x2),
    .io_x3(m_1735_io_x3),
    .io_s(m_1735_io_s),
    .io_cout(m_1735_io_cout)
  );
  Adder m_1736 ( // @[MUL.scala 102:19]
    .io_x1(m_1736_io_x1),
    .io_x2(m_1736_io_x2),
    .io_x3(m_1736_io_x3),
    .io_s(m_1736_io_s),
    .io_cout(m_1736_io_cout)
  );
  Adder m_1737 ( // @[MUL.scala 102:19]
    .io_x1(m_1737_io_x1),
    .io_x2(m_1737_io_x2),
    .io_x3(m_1737_io_x3),
    .io_s(m_1737_io_s),
    .io_cout(m_1737_io_cout)
  );
  Adder m_1738 ( // @[MUL.scala 102:19]
    .io_x1(m_1738_io_x1),
    .io_x2(m_1738_io_x2),
    .io_x3(m_1738_io_x3),
    .io_s(m_1738_io_s),
    .io_cout(m_1738_io_cout)
  );
  Adder m_1739 ( // @[MUL.scala 102:19]
    .io_x1(m_1739_io_x1),
    .io_x2(m_1739_io_x2),
    .io_x3(m_1739_io_x3),
    .io_s(m_1739_io_s),
    .io_cout(m_1739_io_cout)
  );
  Adder m_1740 ( // @[MUL.scala 102:19]
    .io_x1(m_1740_io_x1),
    .io_x2(m_1740_io_x2),
    .io_x3(m_1740_io_x3),
    .io_s(m_1740_io_s),
    .io_cout(m_1740_io_cout)
  );
  Adder m_1741 ( // @[MUL.scala 102:19]
    .io_x1(m_1741_io_x1),
    .io_x2(m_1741_io_x2),
    .io_x3(m_1741_io_x3),
    .io_s(m_1741_io_s),
    .io_cout(m_1741_io_cout)
  );
  Adder m_1742 ( // @[MUL.scala 102:19]
    .io_x1(m_1742_io_x1),
    .io_x2(m_1742_io_x2),
    .io_x3(m_1742_io_x3),
    .io_s(m_1742_io_s),
    .io_cout(m_1742_io_cout)
  );
  Adder m_1743 ( // @[MUL.scala 102:19]
    .io_x1(m_1743_io_x1),
    .io_x2(m_1743_io_x2),
    .io_x3(m_1743_io_x3),
    .io_s(m_1743_io_s),
    .io_cout(m_1743_io_cout)
  );
  Adder m_1744 ( // @[MUL.scala 102:19]
    .io_x1(m_1744_io_x1),
    .io_x2(m_1744_io_x2),
    .io_x3(m_1744_io_x3),
    .io_s(m_1744_io_s),
    .io_cout(m_1744_io_cout)
  );
  Adder m_1745 ( // @[MUL.scala 102:19]
    .io_x1(m_1745_io_x1),
    .io_x2(m_1745_io_x2),
    .io_x3(m_1745_io_x3),
    .io_s(m_1745_io_s),
    .io_cout(m_1745_io_cout)
  );
  Adder m_1746 ( // @[MUL.scala 102:19]
    .io_x1(m_1746_io_x1),
    .io_x2(m_1746_io_x2),
    .io_x3(m_1746_io_x3),
    .io_s(m_1746_io_s),
    .io_cout(m_1746_io_cout)
  );
  Adder m_1747 ( // @[MUL.scala 102:19]
    .io_x1(m_1747_io_x1),
    .io_x2(m_1747_io_x2),
    .io_x3(m_1747_io_x3),
    .io_s(m_1747_io_s),
    .io_cout(m_1747_io_cout)
  );
  Adder m_1748 ( // @[MUL.scala 102:19]
    .io_x1(m_1748_io_x1),
    .io_x2(m_1748_io_x2),
    .io_x3(m_1748_io_x3),
    .io_s(m_1748_io_s),
    .io_cout(m_1748_io_cout)
  );
  Adder m_1749 ( // @[MUL.scala 102:19]
    .io_x1(m_1749_io_x1),
    .io_x2(m_1749_io_x2),
    .io_x3(m_1749_io_x3),
    .io_s(m_1749_io_s),
    .io_cout(m_1749_io_cout)
  );
  Adder m_1750 ( // @[MUL.scala 102:19]
    .io_x1(m_1750_io_x1),
    .io_x2(m_1750_io_x2),
    .io_x3(m_1750_io_x3),
    .io_s(m_1750_io_s),
    .io_cout(m_1750_io_cout)
  );
  Adder m_1751 ( // @[MUL.scala 102:19]
    .io_x1(m_1751_io_x1),
    .io_x2(m_1751_io_x2),
    .io_x3(m_1751_io_x3),
    .io_s(m_1751_io_s),
    .io_cout(m_1751_io_cout)
  );
  Adder m_1752 ( // @[MUL.scala 102:19]
    .io_x1(m_1752_io_x1),
    .io_x2(m_1752_io_x2),
    .io_x3(m_1752_io_x3),
    .io_s(m_1752_io_s),
    .io_cout(m_1752_io_cout)
  );
  Adder m_1753 ( // @[MUL.scala 102:19]
    .io_x1(m_1753_io_x1),
    .io_x2(m_1753_io_x2),
    .io_x3(m_1753_io_x3),
    .io_s(m_1753_io_s),
    .io_cout(m_1753_io_cout)
  );
  Adder m_1754 ( // @[MUL.scala 102:19]
    .io_x1(m_1754_io_x1),
    .io_x2(m_1754_io_x2),
    .io_x3(m_1754_io_x3),
    .io_s(m_1754_io_s),
    .io_cout(m_1754_io_cout)
  );
  Adder m_1755 ( // @[MUL.scala 102:19]
    .io_x1(m_1755_io_x1),
    .io_x2(m_1755_io_x2),
    .io_x3(m_1755_io_x3),
    .io_s(m_1755_io_s),
    .io_cout(m_1755_io_cout)
  );
  Adder m_1756 ( // @[MUL.scala 102:19]
    .io_x1(m_1756_io_x1),
    .io_x2(m_1756_io_x2),
    .io_x3(m_1756_io_x3),
    .io_s(m_1756_io_s),
    .io_cout(m_1756_io_cout)
  );
  Adder m_1757 ( // @[MUL.scala 102:19]
    .io_x1(m_1757_io_x1),
    .io_x2(m_1757_io_x2),
    .io_x3(m_1757_io_x3),
    .io_s(m_1757_io_s),
    .io_cout(m_1757_io_cout)
  );
  Adder m_1758 ( // @[MUL.scala 102:19]
    .io_x1(m_1758_io_x1),
    .io_x2(m_1758_io_x2),
    .io_x3(m_1758_io_x3),
    .io_s(m_1758_io_s),
    .io_cout(m_1758_io_cout)
  );
  Adder m_1759 ( // @[MUL.scala 102:19]
    .io_x1(m_1759_io_x1),
    .io_x2(m_1759_io_x2),
    .io_x3(m_1759_io_x3),
    .io_s(m_1759_io_s),
    .io_cout(m_1759_io_cout)
  );
  Half_Adder m_1760 ( // @[MUL.scala 124:19]
    .io_in_0(m_1760_io_in_0),
    .io_in_1(m_1760_io_in_1),
    .io_out_0(m_1760_io_out_0),
    .io_out_1(m_1760_io_out_1)
  );
  Adder m_1761 ( // @[MUL.scala 102:19]
    .io_x1(m_1761_io_x1),
    .io_x2(m_1761_io_x2),
    .io_x3(m_1761_io_x3),
    .io_s(m_1761_io_s),
    .io_cout(m_1761_io_cout)
  );
  Adder m_1762 ( // @[MUL.scala 102:19]
    .io_x1(m_1762_io_x1),
    .io_x2(m_1762_io_x2),
    .io_x3(m_1762_io_x3),
    .io_s(m_1762_io_s),
    .io_cout(m_1762_io_cout)
  );
  Half_Adder m_1763 ( // @[MUL.scala 124:19]
    .io_in_0(m_1763_io_in_0),
    .io_in_1(m_1763_io_in_1),
    .io_out_0(m_1763_io_out_0),
    .io_out_1(m_1763_io_out_1)
  );
  Adder m_1764 ( // @[MUL.scala 102:19]
    .io_x1(m_1764_io_x1),
    .io_x2(m_1764_io_x2),
    .io_x3(m_1764_io_x3),
    .io_s(m_1764_io_s),
    .io_cout(m_1764_io_cout)
  );
  Adder m_1765 ( // @[MUL.scala 102:19]
    .io_x1(m_1765_io_x1),
    .io_x2(m_1765_io_x2),
    .io_x3(m_1765_io_x3),
    .io_s(m_1765_io_s),
    .io_cout(m_1765_io_cout)
  );
  Half_Adder m_1766 ( // @[MUL.scala 124:19]
    .io_in_0(m_1766_io_in_0),
    .io_in_1(m_1766_io_in_1),
    .io_out_0(m_1766_io_out_0),
    .io_out_1(m_1766_io_out_1)
  );
  Adder m_1767 ( // @[MUL.scala 102:19]
    .io_x1(m_1767_io_x1),
    .io_x2(m_1767_io_x2),
    .io_x3(m_1767_io_x3),
    .io_s(m_1767_io_s),
    .io_cout(m_1767_io_cout)
  );
  Adder m_1768 ( // @[MUL.scala 102:19]
    .io_x1(m_1768_io_x1),
    .io_x2(m_1768_io_x2),
    .io_x3(m_1768_io_x3),
    .io_s(m_1768_io_s),
    .io_cout(m_1768_io_cout)
  );
  Half_Adder m_1769 ( // @[MUL.scala 124:19]
    .io_in_0(m_1769_io_in_0),
    .io_in_1(m_1769_io_in_1),
    .io_out_0(m_1769_io_out_0),
    .io_out_1(m_1769_io_out_1)
  );
  Adder m_1770 ( // @[MUL.scala 102:19]
    .io_x1(m_1770_io_x1),
    .io_x2(m_1770_io_x2),
    .io_x3(m_1770_io_x3),
    .io_s(m_1770_io_s),
    .io_cout(m_1770_io_cout)
  );
  Adder m_1771 ( // @[MUL.scala 102:19]
    .io_x1(m_1771_io_x1),
    .io_x2(m_1771_io_x2),
    .io_x3(m_1771_io_x3),
    .io_s(m_1771_io_s),
    .io_cout(m_1771_io_cout)
  );
  Half_Adder m_1772 ( // @[MUL.scala 124:19]
    .io_in_0(m_1772_io_in_0),
    .io_in_1(m_1772_io_in_1),
    .io_out_0(m_1772_io_out_0),
    .io_out_1(m_1772_io_out_1)
  );
  Adder m_1773 ( // @[MUL.scala 102:19]
    .io_x1(m_1773_io_x1),
    .io_x2(m_1773_io_x2),
    .io_x3(m_1773_io_x3),
    .io_s(m_1773_io_s),
    .io_cout(m_1773_io_cout)
  );
  Adder m_1774 ( // @[MUL.scala 102:19]
    .io_x1(m_1774_io_x1),
    .io_x2(m_1774_io_x2),
    .io_x3(m_1774_io_x3),
    .io_s(m_1774_io_s),
    .io_cout(m_1774_io_cout)
  );
  Half_Adder m_1775 ( // @[MUL.scala 124:19]
    .io_in_0(m_1775_io_in_0),
    .io_in_1(m_1775_io_in_1),
    .io_out_0(m_1775_io_out_0),
    .io_out_1(m_1775_io_out_1)
  );
  Adder m_1776 ( // @[MUL.scala 102:19]
    .io_x1(m_1776_io_x1),
    .io_x2(m_1776_io_x2),
    .io_x3(m_1776_io_x3),
    .io_s(m_1776_io_s),
    .io_cout(m_1776_io_cout)
  );
  Adder m_1777 ( // @[MUL.scala 102:19]
    .io_x1(m_1777_io_x1),
    .io_x2(m_1777_io_x2),
    .io_x3(m_1777_io_x3),
    .io_s(m_1777_io_s),
    .io_cout(m_1777_io_cout)
  );
  Half_Adder m_1778 ( // @[MUL.scala 124:19]
    .io_in_0(m_1778_io_in_0),
    .io_in_1(m_1778_io_in_1),
    .io_out_0(m_1778_io_out_0),
    .io_out_1(m_1778_io_out_1)
  );
  Adder m_1779 ( // @[MUL.scala 102:19]
    .io_x1(m_1779_io_x1),
    .io_x2(m_1779_io_x2),
    .io_x3(m_1779_io_x3),
    .io_s(m_1779_io_s),
    .io_cout(m_1779_io_cout)
  );
  Adder m_1780 ( // @[MUL.scala 102:19]
    .io_x1(m_1780_io_x1),
    .io_x2(m_1780_io_x2),
    .io_x3(m_1780_io_x3),
    .io_s(m_1780_io_s),
    .io_cout(m_1780_io_cout)
  );
  Half_Adder m_1781 ( // @[MUL.scala 124:19]
    .io_in_0(m_1781_io_in_0),
    .io_in_1(m_1781_io_in_1),
    .io_out_0(m_1781_io_out_0),
    .io_out_1(m_1781_io_out_1)
  );
  Adder m_1782 ( // @[MUL.scala 102:19]
    .io_x1(m_1782_io_x1),
    .io_x2(m_1782_io_x2),
    .io_x3(m_1782_io_x3),
    .io_s(m_1782_io_s),
    .io_cout(m_1782_io_cout)
  );
  Adder m_1783 ( // @[MUL.scala 102:19]
    .io_x1(m_1783_io_x1),
    .io_x2(m_1783_io_x2),
    .io_x3(m_1783_io_x3),
    .io_s(m_1783_io_s),
    .io_cout(m_1783_io_cout)
  );
  Adder m_1784 ( // @[MUL.scala 102:19]
    .io_x1(m_1784_io_x1),
    .io_x2(m_1784_io_x2),
    .io_x3(m_1784_io_x3),
    .io_s(m_1784_io_s),
    .io_cout(m_1784_io_cout)
  );
  Adder m_1785 ( // @[MUL.scala 102:19]
    .io_x1(m_1785_io_x1),
    .io_x2(m_1785_io_x2),
    .io_x3(m_1785_io_x3),
    .io_s(m_1785_io_s),
    .io_cout(m_1785_io_cout)
  );
  Adder m_1786 ( // @[MUL.scala 102:19]
    .io_x1(m_1786_io_x1),
    .io_x2(m_1786_io_x2),
    .io_x3(m_1786_io_x3),
    .io_s(m_1786_io_s),
    .io_cout(m_1786_io_cout)
  );
  Adder m_1787 ( // @[MUL.scala 102:19]
    .io_x1(m_1787_io_x1),
    .io_x2(m_1787_io_x2),
    .io_x3(m_1787_io_x3),
    .io_s(m_1787_io_s),
    .io_cout(m_1787_io_cout)
  );
  Adder m_1788 ( // @[MUL.scala 102:19]
    .io_x1(m_1788_io_x1),
    .io_x2(m_1788_io_x2),
    .io_x3(m_1788_io_x3),
    .io_s(m_1788_io_s),
    .io_cout(m_1788_io_cout)
  );
  Adder m_1789 ( // @[MUL.scala 102:19]
    .io_x1(m_1789_io_x1),
    .io_x2(m_1789_io_x2),
    .io_x3(m_1789_io_x3),
    .io_s(m_1789_io_s),
    .io_cout(m_1789_io_cout)
  );
  Adder m_1790 ( // @[MUL.scala 102:19]
    .io_x1(m_1790_io_x1),
    .io_x2(m_1790_io_x2),
    .io_x3(m_1790_io_x3),
    .io_s(m_1790_io_s),
    .io_cout(m_1790_io_cout)
  );
  Adder m_1791 ( // @[MUL.scala 102:19]
    .io_x1(m_1791_io_x1),
    .io_x2(m_1791_io_x2),
    .io_x3(m_1791_io_x3),
    .io_s(m_1791_io_s),
    .io_cout(m_1791_io_cout)
  );
  Adder m_1792 ( // @[MUL.scala 102:19]
    .io_x1(m_1792_io_x1),
    .io_x2(m_1792_io_x2),
    .io_x3(m_1792_io_x3),
    .io_s(m_1792_io_s),
    .io_cout(m_1792_io_cout)
  );
  Adder m_1793 ( // @[MUL.scala 102:19]
    .io_x1(m_1793_io_x1),
    .io_x2(m_1793_io_x2),
    .io_x3(m_1793_io_x3),
    .io_s(m_1793_io_s),
    .io_cout(m_1793_io_cout)
  );
  Adder m_1794 ( // @[MUL.scala 102:19]
    .io_x1(m_1794_io_x1),
    .io_x2(m_1794_io_x2),
    .io_x3(m_1794_io_x3),
    .io_s(m_1794_io_s),
    .io_cout(m_1794_io_cout)
  );
  Adder m_1795 ( // @[MUL.scala 102:19]
    .io_x1(m_1795_io_x1),
    .io_x2(m_1795_io_x2),
    .io_x3(m_1795_io_x3),
    .io_s(m_1795_io_s),
    .io_cout(m_1795_io_cout)
  );
  Adder m_1796 ( // @[MUL.scala 102:19]
    .io_x1(m_1796_io_x1),
    .io_x2(m_1796_io_x2),
    .io_x3(m_1796_io_x3),
    .io_s(m_1796_io_s),
    .io_cout(m_1796_io_cout)
  );
  Adder m_1797 ( // @[MUL.scala 102:19]
    .io_x1(m_1797_io_x1),
    .io_x2(m_1797_io_x2),
    .io_x3(m_1797_io_x3),
    .io_s(m_1797_io_s),
    .io_cout(m_1797_io_cout)
  );
  Adder m_1798 ( // @[MUL.scala 102:19]
    .io_x1(m_1798_io_x1),
    .io_x2(m_1798_io_x2),
    .io_x3(m_1798_io_x3),
    .io_s(m_1798_io_s),
    .io_cout(m_1798_io_cout)
  );
  Adder m_1799 ( // @[MUL.scala 102:19]
    .io_x1(m_1799_io_x1),
    .io_x2(m_1799_io_x2),
    .io_x3(m_1799_io_x3),
    .io_s(m_1799_io_s),
    .io_cout(m_1799_io_cout)
  );
  Adder m_1800 ( // @[MUL.scala 102:19]
    .io_x1(m_1800_io_x1),
    .io_x2(m_1800_io_x2),
    .io_x3(m_1800_io_x3),
    .io_s(m_1800_io_s),
    .io_cout(m_1800_io_cout)
  );
  Adder m_1801 ( // @[MUL.scala 102:19]
    .io_x1(m_1801_io_x1),
    .io_x2(m_1801_io_x2),
    .io_x3(m_1801_io_x3),
    .io_s(m_1801_io_s),
    .io_cout(m_1801_io_cout)
  );
  Adder m_1802 ( // @[MUL.scala 102:19]
    .io_x1(m_1802_io_x1),
    .io_x2(m_1802_io_x2),
    .io_x3(m_1802_io_x3),
    .io_s(m_1802_io_s),
    .io_cout(m_1802_io_cout)
  );
  Adder m_1803 ( // @[MUL.scala 102:19]
    .io_x1(m_1803_io_x1),
    .io_x2(m_1803_io_x2),
    .io_x3(m_1803_io_x3),
    .io_s(m_1803_io_s),
    .io_cout(m_1803_io_cout)
  );
  Adder m_1804 ( // @[MUL.scala 102:19]
    .io_x1(m_1804_io_x1),
    .io_x2(m_1804_io_x2),
    .io_x3(m_1804_io_x3),
    .io_s(m_1804_io_s),
    .io_cout(m_1804_io_cout)
  );
  Adder m_1805 ( // @[MUL.scala 102:19]
    .io_x1(m_1805_io_x1),
    .io_x2(m_1805_io_x2),
    .io_x3(m_1805_io_x3),
    .io_s(m_1805_io_s),
    .io_cout(m_1805_io_cout)
  );
  Adder m_1806 ( // @[MUL.scala 102:19]
    .io_x1(m_1806_io_x1),
    .io_x2(m_1806_io_x2),
    .io_x3(m_1806_io_x3),
    .io_s(m_1806_io_s),
    .io_cout(m_1806_io_cout)
  );
  Adder m_1807 ( // @[MUL.scala 102:19]
    .io_x1(m_1807_io_x1),
    .io_x2(m_1807_io_x2),
    .io_x3(m_1807_io_x3),
    .io_s(m_1807_io_s),
    .io_cout(m_1807_io_cout)
  );
  Adder m_1808 ( // @[MUL.scala 102:19]
    .io_x1(m_1808_io_x1),
    .io_x2(m_1808_io_x2),
    .io_x3(m_1808_io_x3),
    .io_s(m_1808_io_s),
    .io_cout(m_1808_io_cout)
  );
  Adder m_1809 ( // @[MUL.scala 102:19]
    .io_x1(m_1809_io_x1),
    .io_x2(m_1809_io_x2),
    .io_x3(m_1809_io_x3),
    .io_s(m_1809_io_s),
    .io_cout(m_1809_io_cout)
  );
  Adder m_1810 ( // @[MUL.scala 102:19]
    .io_x1(m_1810_io_x1),
    .io_x2(m_1810_io_x2),
    .io_x3(m_1810_io_x3),
    .io_s(m_1810_io_s),
    .io_cout(m_1810_io_cout)
  );
  Adder m_1811 ( // @[MUL.scala 102:19]
    .io_x1(m_1811_io_x1),
    .io_x2(m_1811_io_x2),
    .io_x3(m_1811_io_x3),
    .io_s(m_1811_io_s),
    .io_cout(m_1811_io_cout)
  );
  Adder m_1812 ( // @[MUL.scala 102:19]
    .io_x1(m_1812_io_x1),
    .io_x2(m_1812_io_x2),
    .io_x3(m_1812_io_x3),
    .io_s(m_1812_io_s),
    .io_cout(m_1812_io_cout)
  );
  Adder m_1813 ( // @[MUL.scala 102:19]
    .io_x1(m_1813_io_x1),
    .io_x2(m_1813_io_x2),
    .io_x3(m_1813_io_x3),
    .io_s(m_1813_io_s),
    .io_cout(m_1813_io_cout)
  );
  Adder m_1814 ( // @[MUL.scala 102:19]
    .io_x1(m_1814_io_x1),
    .io_x2(m_1814_io_x2),
    .io_x3(m_1814_io_x3),
    .io_s(m_1814_io_s),
    .io_cout(m_1814_io_cout)
  );
  Adder m_1815 ( // @[MUL.scala 102:19]
    .io_x1(m_1815_io_x1),
    .io_x2(m_1815_io_x2),
    .io_x3(m_1815_io_x3),
    .io_s(m_1815_io_s),
    .io_cout(m_1815_io_cout)
  );
  Adder m_1816 ( // @[MUL.scala 102:19]
    .io_x1(m_1816_io_x1),
    .io_x2(m_1816_io_x2),
    .io_x3(m_1816_io_x3),
    .io_s(m_1816_io_s),
    .io_cout(m_1816_io_cout)
  );
  Adder m_1817 ( // @[MUL.scala 102:19]
    .io_x1(m_1817_io_x1),
    .io_x2(m_1817_io_x2),
    .io_x3(m_1817_io_x3),
    .io_s(m_1817_io_s),
    .io_cout(m_1817_io_cout)
  );
  Adder m_1818 ( // @[MUL.scala 102:19]
    .io_x1(m_1818_io_x1),
    .io_x2(m_1818_io_x2),
    .io_x3(m_1818_io_x3),
    .io_s(m_1818_io_s),
    .io_cout(m_1818_io_cout)
  );
  Adder m_1819 ( // @[MUL.scala 102:19]
    .io_x1(m_1819_io_x1),
    .io_x2(m_1819_io_x2),
    .io_x3(m_1819_io_x3),
    .io_s(m_1819_io_s),
    .io_cout(m_1819_io_cout)
  );
  Adder m_1820 ( // @[MUL.scala 102:19]
    .io_x1(m_1820_io_x1),
    .io_x2(m_1820_io_x2),
    .io_x3(m_1820_io_x3),
    .io_s(m_1820_io_s),
    .io_cout(m_1820_io_cout)
  );
  Adder m_1821 ( // @[MUL.scala 102:19]
    .io_x1(m_1821_io_x1),
    .io_x2(m_1821_io_x2),
    .io_x3(m_1821_io_x3),
    .io_s(m_1821_io_s),
    .io_cout(m_1821_io_cout)
  );
  Adder m_1822 ( // @[MUL.scala 102:19]
    .io_x1(m_1822_io_x1),
    .io_x2(m_1822_io_x2),
    .io_x3(m_1822_io_x3),
    .io_s(m_1822_io_s),
    .io_cout(m_1822_io_cout)
  );
  Adder m_1823 ( // @[MUL.scala 102:19]
    .io_x1(m_1823_io_x1),
    .io_x2(m_1823_io_x2),
    .io_x3(m_1823_io_x3),
    .io_s(m_1823_io_s),
    .io_cout(m_1823_io_cout)
  );
  Adder m_1824 ( // @[MUL.scala 102:19]
    .io_x1(m_1824_io_x1),
    .io_x2(m_1824_io_x2),
    .io_x3(m_1824_io_x3),
    .io_s(m_1824_io_s),
    .io_cout(m_1824_io_cout)
  );
  Adder m_1825 ( // @[MUL.scala 102:19]
    .io_x1(m_1825_io_x1),
    .io_x2(m_1825_io_x2),
    .io_x3(m_1825_io_x3),
    .io_s(m_1825_io_s),
    .io_cout(m_1825_io_cout)
  );
  Adder m_1826 ( // @[MUL.scala 102:19]
    .io_x1(m_1826_io_x1),
    .io_x2(m_1826_io_x2),
    .io_x3(m_1826_io_x3),
    .io_s(m_1826_io_s),
    .io_cout(m_1826_io_cout)
  );
  Adder m_1827 ( // @[MUL.scala 102:19]
    .io_x1(m_1827_io_x1),
    .io_x2(m_1827_io_x2),
    .io_x3(m_1827_io_x3),
    .io_s(m_1827_io_s),
    .io_cout(m_1827_io_cout)
  );
  Adder m_1828 ( // @[MUL.scala 102:19]
    .io_x1(m_1828_io_x1),
    .io_x2(m_1828_io_x2),
    .io_x3(m_1828_io_x3),
    .io_s(m_1828_io_s),
    .io_cout(m_1828_io_cout)
  );
  Adder m_1829 ( // @[MUL.scala 102:19]
    .io_x1(m_1829_io_x1),
    .io_x2(m_1829_io_x2),
    .io_x3(m_1829_io_x3),
    .io_s(m_1829_io_s),
    .io_cout(m_1829_io_cout)
  );
  Adder m_1830 ( // @[MUL.scala 102:19]
    .io_x1(m_1830_io_x1),
    .io_x2(m_1830_io_x2),
    .io_x3(m_1830_io_x3),
    .io_s(m_1830_io_s),
    .io_cout(m_1830_io_cout)
  );
  Adder m_1831 ( // @[MUL.scala 102:19]
    .io_x1(m_1831_io_x1),
    .io_x2(m_1831_io_x2),
    .io_x3(m_1831_io_x3),
    .io_s(m_1831_io_s),
    .io_cout(m_1831_io_cout)
  );
  Adder m_1832 ( // @[MUL.scala 102:19]
    .io_x1(m_1832_io_x1),
    .io_x2(m_1832_io_x2),
    .io_x3(m_1832_io_x3),
    .io_s(m_1832_io_s),
    .io_cout(m_1832_io_cout)
  );
  Adder m_1833 ( // @[MUL.scala 102:19]
    .io_x1(m_1833_io_x1),
    .io_x2(m_1833_io_x2),
    .io_x3(m_1833_io_x3),
    .io_s(m_1833_io_s),
    .io_cout(m_1833_io_cout)
  );
  Adder m_1834 ( // @[MUL.scala 102:19]
    .io_x1(m_1834_io_x1),
    .io_x2(m_1834_io_x2),
    .io_x3(m_1834_io_x3),
    .io_s(m_1834_io_s),
    .io_cout(m_1834_io_cout)
  );
  Adder m_1835 ( // @[MUL.scala 102:19]
    .io_x1(m_1835_io_x1),
    .io_x2(m_1835_io_x2),
    .io_x3(m_1835_io_x3),
    .io_s(m_1835_io_s),
    .io_cout(m_1835_io_cout)
  );
  Adder m_1836 ( // @[MUL.scala 102:19]
    .io_x1(m_1836_io_x1),
    .io_x2(m_1836_io_x2),
    .io_x3(m_1836_io_x3),
    .io_s(m_1836_io_s),
    .io_cout(m_1836_io_cout)
  );
  Adder m_1837 ( // @[MUL.scala 102:19]
    .io_x1(m_1837_io_x1),
    .io_x2(m_1837_io_x2),
    .io_x3(m_1837_io_x3),
    .io_s(m_1837_io_s),
    .io_cout(m_1837_io_cout)
  );
  Adder m_1838 ( // @[MUL.scala 102:19]
    .io_x1(m_1838_io_x1),
    .io_x2(m_1838_io_x2),
    .io_x3(m_1838_io_x3),
    .io_s(m_1838_io_s),
    .io_cout(m_1838_io_cout)
  );
  Adder m_1839 ( // @[MUL.scala 102:19]
    .io_x1(m_1839_io_x1),
    .io_x2(m_1839_io_x2),
    .io_x3(m_1839_io_x3),
    .io_s(m_1839_io_s),
    .io_cout(m_1839_io_cout)
  );
  Adder m_1840 ( // @[MUL.scala 102:19]
    .io_x1(m_1840_io_x1),
    .io_x2(m_1840_io_x2),
    .io_x3(m_1840_io_x3),
    .io_s(m_1840_io_s),
    .io_cout(m_1840_io_cout)
  );
  Adder m_1841 ( // @[MUL.scala 102:19]
    .io_x1(m_1841_io_x1),
    .io_x2(m_1841_io_x2),
    .io_x3(m_1841_io_x3),
    .io_s(m_1841_io_s),
    .io_cout(m_1841_io_cout)
  );
  Adder m_1842 ( // @[MUL.scala 102:19]
    .io_x1(m_1842_io_x1),
    .io_x2(m_1842_io_x2),
    .io_x3(m_1842_io_x3),
    .io_s(m_1842_io_s),
    .io_cout(m_1842_io_cout)
  );
  Adder m_1843 ( // @[MUL.scala 102:19]
    .io_x1(m_1843_io_x1),
    .io_x2(m_1843_io_x2),
    .io_x3(m_1843_io_x3),
    .io_s(m_1843_io_s),
    .io_cout(m_1843_io_cout)
  );
  Adder m_1844 ( // @[MUL.scala 102:19]
    .io_x1(m_1844_io_x1),
    .io_x2(m_1844_io_x2),
    .io_x3(m_1844_io_x3),
    .io_s(m_1844_io_s),
    .io_cout(m_1844_io_cout)
  );
  Adder m_1845 ( // @[MUL.scala 102:19]
    .io_x1(m_1845_io_x1),
    .io_x2(m_1845_io_x2),
    .io_x3(m_1845_io_x3),
    .io_s(m_1845_io_s),
    .io_cout(m_1845_io_cout)
  );
  Adder m_1846 ( // @[MUL.scala 102:19]
    .io_x1(m_1846_io_x1),
    .io_x2(m_1846_io_x2),
    .io_x3(m_1846_io_x3),
    .io_s(m_1846_io_s),
    .io_cout(m_1846_io_cout)
  );
  Adder m_1847 ( // @[MUL.scala 102:19]
    .io_x1(m_1847_io_x1),
    .io_x2(m_1847_io_x2),
    .io_x3(m_1847_io_x3),
    .io_s(m_1847_io_s),
    .io_cout(m_1847_io_cout)
  );
  Adder m_1848 ( // @[MUL.scala 102:19]
    .io_x1(m_1848_io_x1),
    .io_x2(m_1848_io_x2),
    .io_x3(m_1848_io_x3),
    .io_s(m_1848_io_s),
    .io_cout(m_1848_io_cout)
  );
  Adder m_1849 ( // @[MUL.scala 102:19]
    .io_x1(m_1849_io_x1),
    .io_x2(m_1849_io_x2),
    .io_x3(m_1849_io_x3),
    .io_s(m_1849_io_s),
    .io_cout(m_1849_io_cout)
  );
  Adder m_1850 ( // @[MUL.scala 102:19]
    .io_x1(m_1850_io_x1),
    .io_x2(m_1850_io_x2),
    .io_x3(m_1850_io_x3),
    .io_s(m_1850_io_s),
    .io_cout(m_1850_io_cout)
  );
  Adder m_1851 ( // @[MUL.scala 102:19]
    .io_x1(m_1851_io_x1),
    .io_x2(m_1851_io_x2),
    .io_x3(m_1851_io_x3),
    .io_s(m_1851_io_s),
    .io_cout(m_1851_io_cout)
  );
  Adder m_1852 ( // @[MUL.scala 102:19]
    .io_x1(m_1852_io_x1),
    .io_x2(m_1852_io_x2),
    .io_x3(m_1852_io_x3),
    .io_s(m_1852_io_s),
    .io_cout(m_1852_io_cout)
  );
  Adder m_1853 ( // @[MUL.scala 102:19]
    .io_x1(m_1853_io_x1),
    .io_x2(m_1853_io_x2),
    .io_x3(m_1853_io_x3),
    .io_s(m_1853_io_s),
    .io_cout(m_1853_io_cout)
  );
  Adder m_1854 ( // @[MUL.scala 102:19]
    .io_x1(m_1854_io_x1),
    .io_x2(m_1854_io_x2),
    .io_x3(m_1854_io_x3),
    .io_s(m_1854_io_s),
    .io_cout(m_1854_io_cout)
  );
  Adder m_1855 ( // @[MUL.scala 102:19]
    .io_x1(m_1855_io_x1),
    .io_x2(m_1855_io_x2),
    .io_x3(m_1855_io_x3),
    .io_s(m_1855_io_s),
    .io_cout(m_1855_io_cout)
  );
  Adder m_1856 ( // @[MUL.scala 102:19]
    .io_x1(m_1856_io_x1),
    .io_x2(m_1856_io_x2),
    .io_x3(m_1856_io_x3),
    .io_s(m_1856_io_s),
    .io_cout(m_1856_io_cout)
  );
  Adder m_1857 ( // @[MUL.scala 102:19]
    .io_x1(m_1857_io_x1),
    .io_x2(m_1857_io_x2),
    .io_x3(m_1857_io_x3),
    .io_s(m_1857_io_s),
    .io_cout(m_1857_io_cout)
  );
  Adder m_1858 ( // @[MUL.scala 102:19]
    .io_x1(m_1858_io_x1),
    .io_x2(m_1858_io_x2),
    .io_x3(m_1858_io_x3),
    .io_s(m_1858_io_s),
    .io_cout(m_1858_io_cout)
  );
  Adder m_1859 ( // @[MUL.scala 102:19]
    .io_x1(m_1859_io_x1),
    .io_x2(m_1859_io_x2),
    .io_x3(m_1859_io_x3),
    .io_s(m_1859_io_s),
    .io_cout(m_1859_io_cout)
  );
  Adder m_1860 ( // @[MUL.scala 102:19]
    .io_x1(m_1860_io_x1),
    .io_x2(m_1860_io_x2),
    .io_x3(m_1860_io_x3),
    .io_s(m_1860_io_s),
    .io_cout(m_1860_io_cout)
  );
  Adder m_1861 ( // @[MUL.scala 102:19]
    .io_x1(m_1861_io_x1),
    .io_x2(m_1861_io_x2),
    .io_x3(m_1861_io_x3),
    .io_s(m_1861_io_s),
    .io_cout(m_1861_io_cout)
  );
  Adder m_1862 ( // @[MUL.scala 102:19]
    .io_x1(m_1862_io_x1),
    .io_x2(m_1862_io_x2),
    .io_x3(m_1862_io_x3),
    .io_s(m_1862_io_s),
    .io_cout(m_1862_io_cout)
  );
  Adder m_1863 ( // @[MUL.scala 102:19]
    .io_x1(m_1863_io_x1),
    .io_x2(m_1863_io_x2),
    .io_x3(m_1863_io_x3),
    .io_s(m_1863_io_s),
    .io_cout(m_1863_io_cout)
  );
  Adder m_1864 ( // @[MUL.scala 102:19]
    .io_x1(m_1864_io_x1),
    .io_x2(m_1864_io_x2),
    .io_x3(m_1864_io_x3),
    .io_s(m_1864_io_s),
    .io_cout(m_1864_io_cout)
  );
  Half_Adder m_1865 ( // @[MUL.scala 124:19]
    .io_in_0(m_1865_io_in_0),
    .io_in_1(m_1865_io_in_1),
    .io_out_0(m_1865_io_out_0),
    .io_out_1(m_1865_io_out_1)
  );
  Adder m_1866 ( // @[MUL.scala 102:19]
    .io_x1(m_1866_io_x1),
    .io_x2(m_1866_io_x2),
    .io_x3(m_1866_io_x3),
    .io_s(m_1866_io_s),
    .io_cout(m_1866_io_cout)
  );
  Adder m_1867 ( // @[MUL.scala 102:19]
    .io_x1(m_1867_io_x1),
    .io_x2(m_1867_io_x2),
    .io_x3(m_1867_io_x3),
    .io_s(m_1867_io_s),
    .io_cout(m_1867_io_cout)
  );
  Half_Adder m_1868 ( // @[MUL.scala 124:19]
    .io_in_0(m_1868_io_in_0),
    .io_in_1(m_1868_io_in_1),
    .io_out_0(m_1868_io_out_0),
    .io_out_1(m_1868_io_out_1)
  );
  Adder m_1869 ( // @[MUL.scala 102:19]
    .io_x1(m_1869_io_x1),
    .io_x2(m_1869_io_x2),
    .io_x3(m_1869_io_x3),
    .io_s(m_1869_io_s),
    .io_cout(m_1869_io_cout)
  );
  Adder m_1870 ( // @[MUL.scala 102:19]
    .io_x1(m_1870_io_x1),
    .io_x2(m_1870_io_x2),
    .io_x3(m_1870_io_x3),
    .io_s(m_1870_io_s),
    .io_cout(m_1870_io_cout)
  );
  Half_Adder m_1871 ( // @[MUL.scala 124:19]
    .io_in_0(m_1871_io_in_0),
    .io_in_1(m_1871_io_in_1),
    .io_out_0(m_1871_io_out_0),
    .io_out_1(m_1871_io_out_1)
  );
  Adder m_1872 ( // @[MUL.scala 102:19]
    .io_x1(m_1872_io_x1),
    .io_x2(m_1872_io_x2),
    .io_x3(m_1872_io_x3),
    .io_s(m_1872_io_s),
    .io_cout(m_1872_io_cout)
  );
  Adder m_1873 ( // @[MUL.scala 102:19]
    .io_x1(m_1873_io_x1),
    .io_x2(m_1873_io_x2),
    .io_x3(m_1873_io_x3),
    .io_s(m_1873_io_s),
    .io_cout(m_1873_io_cout)
  );
  Half_Adder m_1874 ( // @[MUL.scala 124:19]
    .io_in_0(m_1874_io_in_0),
    .io_in_1(m_1874_io_in_1),
    .io_out_0(m_1874_io_out_0),
    .io_out_1(m_1874_io_out_1)
  );
  Adder m_1875 ( // @[MUL.scala 102:19]
    .io_x1(m_1875_io_x1),
    .io_x2(m_1875_io_x2),
    .io_x3(m_1875_io_x3),
    .io_s(m_1875_io_s),
    .io_cout(m_1875_io_cout)
  );
  Adder m_1876 ( // @[MUL.scala 102:19]
    .io_x1(m_1876_io_x1),
    .io_x2(m_1876_io_x2),
    .io_x3(m_1876_io_x3),
    .io_s(m_1876_io_s),
    .io_cout(m_1876_io_cout)
  );
  Half_Adder m_1877 ( // @[MUL.scala 124:19]
    .io_in_0(m_1877_io_in_0),
    .io_in_1(m_1877_io_in_1),
    .io_out_0(m_1877_io_out_0),
    .io_out_1(m_1877_io_out_1)
  );
  Adder m_1878 ( // @[MUL.scala 102:19]
    .io_x1(m_1878_io_x1),
    .io_x2(m_1878_io_x2),
    .io_x3(m_1878_io_x3),
    .io_s(m_1878_io_s),
    .io_cout(m_1878_io_cout)
  );
  Adder m_1879 ( // @[MUL.scala 102:19]
    .io_x1(m_1879_io_x1),
    .io_x2(m_1879_io_x2),
    .io_x3(m_1879_io_x3),
    .io_s(m_1879_io_s),
    .io_cout(m_1879_io_cout)
  );
  Half_Adder m_1880 ( // @[MUL.scala 124:19]
    .io_in_0(m_1880_io_in_0),
    .io_in_1(m_1880_io_in_1),
    .io_out_0(m_1880_io_out_0),
    .io_out_1(m_1880_io_out_1)
  );
  Adder m_1881 ( // @[MUL.scala 102:19]
    .io_x1(m_1881_io_x1),
    .io_x2(m_1881_io_x2),
    .io_x3(m_1881_io_x3),
    .io_s(m_1881_io_s),
    .io_cout(m_1881_io_cout)
  );
  Adder m_1882 ( // @[MUL.scala 102:19]
    .io_x1(m_1882_io_x1),
    .io_x2(m_1882_io_x2),
    .io_x3(m_1882_io_x3),
    .io_s(m_1882_io_s),
    .io_cout(m_1882_io_cout)
  );
  Half_Adder m_1883 ( // @[MUL.scala 124:19]
    .io_in_0(m_1883_io_in_0),
    .io_in_1(m_1883_io_in_1),
    .io_out_0(m_1883_io_out_0),
    .io_out_1(m_1883_io_out_1)
  );
  Adder m_1884 ( // @[MUL.scala 102:19]
    .io_x1(m_1884_io_x1),
    .io_x2(m_1884_io_x2),
    .io_x3(m_1884_io_x3),
    .io_s(m_1884_io_s),
    .io_cout(m_1884_io_cout)
  );
  Adder m_1885 ( // @[MUL.scala 102:19]
    .io_x1(m_1885_io_x1),
    .io_x2(m_1885_io_x2),
    .io_x3(m_1885_io_x3),
    .io_s(m_1885_io_s),
    .io_cout(m_1885_io_cout)
  );
  Half_Adder m_1886 ( // @[MUL.scala 124:19]
    .io_in_0(m_1886_io_in_0),
    .io_in_1(m_1886_io_in_1),
    .io_out_0(m_1886_io_out_0),
    .io_out_1(m_1886_io_out_1)
  );
  Adder m_1887 ( // @[MUL.scala 102:19]
    .io_x1(m_1887_io_x1),
    .io_x2(m_1887_io_x2),
    .io_x3(m_1887_io_x3),
    .io_s(m_1887_io_s),
    .io_cout(m_1887_io_cout)
  );
  Adder m_1888 ( // @[MUL.scala 102:19]
    .io_x1(m_1888_io_x1),
    .io_x2(m_1888_io_x2),
    .io_x3(m_1888_io_x3),
    .io_s(m_1888_io_s),
    .io_cout(m_1888_io_cout)
  );
  Half_Adder m_1889 ( // @[MUL.scala 124:19]
    .io_in_0(m_1889_io_in_0),
    .io_in_1(m_1889_io_in_1),
    .io_out_0(m_1889_io_out_0),
    .io_out_1(m_1889_io_out_1)
  );
  Adder m_1890 ( // @[MUL.scala 102:19]
    .io_x1(m_1890_io_x1),
    .io_x2(m_1890_io_x2),
    .io_x3(m_1890_io_x3),
    .io_s(m_1890_io_s),
    .io_cout(m_1890_io_cout)
  );
  Adder m_1891 ( // @[MUL.scala 102:19]
    .io_x1(m_1891_io_x1),
    .io_x2(m_1891_io_x2),
    .io_x3(m_1891_io_x3),
    .io_s(m_1891_io_s),
    .io_cout(m_1891_io_cout)
  );
  Half_Adder m_1892 ( // @[MUL.scala 124:19]
    .io_in_0(m_1892_io_in_0),
    .io_in_1(m_1892_io_in_1),
    .io_out_0(m_1892_io_out_0),
    .io_out_1(m_1892_io_out_1)
  );
  Adder m_1893 ( // @[MUL.scala 102:19]
    .io_x1(m_1893_io_x1),
    .io_x2(m_1893_io_x2),
    .io_x3(m_1893_io_x3),
    .io_s(m_1893_io_s),
    .io_cout(m_1893_io_cout)
  );
  Adder m_1894 ( // @[MUL.scala 102:19]
    .io_x1(m_1894_io_x1),
    .io_x2(m_1894_io_x2),
    .io_x3(m_1894_io_x3),
    .io_s(m_1894_io_s),
    .io_cout(m_1894_io_cout)
  );
  Half_Adder m_1895 ( // @[MUL.scala 124:19]
    .io_in_0(m_1895_io_in_0),
    .io_in_1(m_1895_io_in_1),
    .io_out_0(m_1895_io_out_0),
    .io_out_1(m_1895_io_out_1)
  );
  Adder m_1896 ( // @[MUL.scala 102:19]
    .io_x1(m_1896_io_x1),
    .io_x2(m_1896_io_x2),
    .io_x3(m_1896_io_x3),
    .io_s(m_1896_io_s),
    .io_cout(m_1896_io_cout)
  );
  Adder m_1897 ( // @[MUL.scala 102:19]
    .io_x1(m_1897_io_x1),
    .io_x2(m_1897_io_x2),
    .io_x3(m_1897_io_x3),
    .io_s(m_1897_io_s),
    .io_cout(m_1897_io_cout)
  );
  Adder m_1898 ( // @[MUL.scala 102:19]
    .io_x1(m_1898_io_x1),
    .io_x2(m_1898_io_x2),
    .io_x3(m_1898_io_x3),
    .io_s(m_1898_io_s),
    .io_cout(m_1898_io_cout)
  );
  Adder m_1899 ( // @[MUL.scala 102:19]
    .io_x1(m_1899_io_x1),
    .io_x2(m_1899_io_x2),
    .io_x3(m_1899_io_x3),
    .io_s(m_1899_io_s),
    .io_cout(m_1899_io_cout)
  );
  Adder m_1900 ( // @[MUL.scala 102:19]
    .io_x1(m_1900_io_x1),
    .io_x2(m_1900_io_x2),
    .io_x3(m_1900_io_x3),
    .io_s(m_1900_io_s),
    .io_cout(m_1900_io_cout)
  );
  Adder m_1901 ( // @[MUL.scala 102:19]
    .io_x1(m_1901_io_x1),
    .io_x2(m_1901_io_x2),
    .io_x3(m_1901_io_x3),
    .io_s(m_1901_io_s),
    .io_cout(m_1901_io_cout)
  );
  Adder m_1902 ( // @[MUL.scala 102:19]
    .io_x1(m_1902_io_x1),
    .io_x2(m_1902_io_x2),
    .io_x3(m_1902_io_x3),
    .io_s(m_1902_io_s),
    .io_cout(m_1902_io_cout)
  );
  Adder m_1903 ( // @[MUL.scala 102:19]
    .io_x1(m_1903_io_x1),
    .io_x2(m_1903_io_x2),
    .io_x3(m_1903_io_x3),
    .io_s(m_1903_io_s),
    .io_cout(m_1903_io_cout)
  );
  Adder m_1904 ( // @[MUL.scala 102:19]
    .io_x1(m_1904_io_x1),
    .io_x2(m_1904_io_x2),
    .io_x3(m_1904_io_x3),
    .io_s(m_1904_io_s),
    .io_cout(m_1904_io_cout)
  );
  Adder m_1905 ( // @[MUL.scala 102:19]
    .io_x1(m_1905_io_x1),
    .io_x2(m_1905_io_x2),
    .io_x3(m_1905_io_x3),
    .io_s(m_1905_io_s),
    .io_cout(m_1905_io_cout)
  );
  Adder m_1906 ( // @[MUL.scala 102:19]
    .io_x1(m_1906_io_x1),
    .io_x2(m_1906_io_x2),
    .io_x3(m_1906_io_x3),
    .io_s(m_1906_io_s),
    .io_cout(m_1906_io_cout)
  );
  Adder m_1907 ( // @[MUL.scala 102:19]
    .io_x1(m_1907_io_x1),
    .io_x2(m_1907_io_x2),
    .io_x3(m_1907_io_x3),
    .io_s(m_1907_io_s),
    .io_cout(m_1907_io_cout)
  );
  Adder m_1908 ( // @[MUL.scala 102:19]
    .io_x1(m_1908_io_x1),
    .io_x2(m_1908_io_x2),
    .io_x3(m_1908_io_x3),
    .io_s(m_1908_io_s),
    .io_cout(m_1908_io_cout)
  );
  Adder m_1909 ( // @[MUL.scala 102:19]
    .io_x1(m_1909_io_x1),
    .io_x2(m_1909_io_x2),
    .io_x3(m_1909_io_x3),
    .io_s(m_1909_io_s),
    .io_cout(m_1909_io_cout)
  );
  Adder m_1910 ( // @[MUL.scala 102:19]
    .io_x1(m_1910_io_x1),
    .io_x2(m_1910_io_x2),
    .io_x3(m_1910_io_x3),
    .io_s(m_1910_io_s),
    .io_cout(m_1910_io_cout)
  );
  Adder m_1911 ( // @[MUL.scala 102:19]
    .io_x1(m_1911_io_x1),
    .io_x2(m_1911_io_x2),
    .io_x3(m_1911_io_x3),
    .io_s(m_1911_io_s),
    .io_cout(m_1911_io_cout)
  );
  Adder m_1912 ( // @[MUL.scala 102:19]
    .io_x1(m_1912_io_x1),
    .io_x2(m_1912_io_x2),
    .io_x3(m_1912_io_x3),
    .io_s(m_1912_io_s),
    .io_cout(m_1912_io_cout)
  );
  Adder m_1913 ( // @[MUL.scala 102:19]
    .io_x1(m_1913_io_x1),
    .io_x2(m_1913_io_x2),
    .io_x3(m_1913_io_x3),
    .io_s(m_1913_io_s),
    .io_cout(m_1913_io_cout)
  );
  Adder m_1914 ( // @[MUL.scala 102:19]
    .io_x1(m_1914_io_x1),
    .io_x2(m_1914_io_x2),
    .io_x3(m_1914_io_x3),
    .io_s(m_1914_io_s),
    .io_cout(m_1914_io_cout)
  );
  Adder m_1915 ( // @[MUL.scala 102:19]
    .io_x1(m_1915_io_x1),
    .io_x2(m_1915_io_x2),
    .io_x3(m_1915_io_x3),
    .io_s(m_1915_io_s),
    .io_cout(m_1915_io_cout)
  );
  Adder m_1916 ( // @[MUL.scala 102:19]
    .io_x1(m_1916_io_x1),
    .io_x2(m_1916_io_x2),
    .io_x3(m_1916_io_x3),
    .io_s(m_1916_io_s),
    .io_cout(m_1916_io_cout)
  );
  Adder m_1917 ( // @[MUL.scala 102:19]
    .io_x1(m_1917_io_x1),
    .io_x2(m_1917_io_x2),
    .io_x3(m_1917_io_x3),
    .io_s(m_1917_io_s),
    .io_cout(m_1917_io_cout)
  );
  Adder m_1918 ( // @[MUL.scala 102:19]
    .io_x1(m_1918_io_x1),
    .io_x2(m_1918_io_x2),
    .io_x3(m_1918_io_x3),
    .io_s(m_1918_io_s),
    .io_cout(m_1918_io_cout)
  );
  Adder m_1919 ( // @[MUL.scala 102:19]
    .io_x1(m_1919_io_x1),
    .io_x2(m_1919_io_x2),
    .io_x3(m_1919_io_x3),
    .io_s(m_1919_io_s),
    .io_cout(m_1919_io_cout)
  );
  Adder m_1920 ( // @[MUL.scala 102:19]
    .io_x1(m_1920_io_x1),
    .io_x2(m_1920_io_x2),
    .io_x3(m_1920_io_x3),
    .io_s(m_1920_io_s),
    .io_cout(m_1920_io_cout)
  );
  Adder m_1921 ( // @[MUL.scala 102:19]
    .io_x1(m_1921_io_x1),
    .io_x2(m_1921_io_x2),
    .io_x3(m_1921_io_x3),
    .io_s(m_1921_io_s),
    .io_cout(m_1921_io_cout)
  );
  Adder m_1922 ( // @[MUL.scala 102:19]
    .io_x1(m_1922_io_x1),
    .io_x2(m_1922_io_x2),
    .io_x3(m_1922_io_x3),
    .io_s(m_1922_io_s),
    .io_cout(m_1922_io_cout)
  );
  Adder m_1923 ( // @[MUL.scala 102:19]
    .io_x1(m_1923_io_x1),
    .io_x2(m_1923_io_x2),
    .io_x3(m_1923_io_x3),
    .io_s(m_1923_io_s),
    .io_cout(m_1923_io_cout)
  );
  Adder m_1924 ( // @[MUL.scala 102:19]
    .io_x1(m_1924_io_x1),
    .io_x2(m_1924_io_x2),
    .io_x3(m_1924_io_x3),
    .io_s(m_1924_io_s),
    .io_cout(m_1924_io_cout)
  );
  Half_Adder m_1925 ( // @[MUL.scala 124:19]
    .io_in_0(m_1925_io_in_0),
    .io_in_1(m_1925_io_in_1),
    .io_out_0(m_1925_io_out_0),
    .io_out_1(m_1925_io_out_1)
  );
  Adder m_1926 ( // @[MUL.scala 102:19]
    .io_x1(m_1926_io_x1),
    .io_x2(m_1926_io_x2),
    .io_x3(m_1926_io_x3),
    .io_s(m_1926_io_s),
    .io_cout(m_1926_io_cout)
  );
  Half_Adder m_1927 ( // @[MUL.scala 124:19]
    .io_in_0(m_1927_io_in_0),
    .io_in_1(m_1927_io_in_1),
    .io_out_0(m_1927_io_out_0),
    .io_out_1(m_1927_io_out_1)
  );
  Adder m_1928 ( // @[MUL.scala 102:19]
    .io_x1(m_1928_io_x1),
    .io_x2(m_1928_io_x2),
    .io_x3(m_1928_io_x3),
    .io_s(m_1928_io_s),
    .io_cout(m_1928_io_cout)
  );
  Half_Adder m_1929 ( // @[MUL.scala 124:19]
    .io_in_0(m_1929_io_in_0),
    .io_in_1(m_1929_io_in_1),
    .io_out_0(m_1929_io_out_0),
    .io_out_1(m_1929_io_out_1)
  );
  Adder m_1930 ( // @[MUL.scala 102:19]
    .io_x1(m_1930_io_x1),
    .io_x2(m_1930_io_x2),
    .io_x3(m_1930_io_x3),
    .io_s(m_1930_io_s),
    .io_cout(m_1930_io_cout)
  );
  Adder m_1931 ( // @[MUL.scala 102:19]
    .io_x1(m_1931_io_x1),
    .io_x2(m_1931_io_x2),
    .io_x3(m_1931_io_x3),
    .io_s(m_1931_io_s),
    .io_cout(m_1931_io_cout)
  );
  Adder m_1932 ( // @[MUL.scala 102:19]
    .io_x1(m_1932_io_x1),
    .io_x2(m_1932_io_x2),
    .io_x3(m_1932_io_x3),
    .io_s(m_1932_io_s),
    .io_cout(m_1932_io_cout)
  );
  Adder m_1933 ( // @[MUL.scala 102:19]
    .io_x1(m_1933_io_x1),
    .io_x2(m_1933_io_x2),
    .io_x3(m_1933_io_x3),
    .io_s(m_1933_io_s),
    .io_cout(m_1933_io_cout)
  );
  Adder m_1934 ( // @[MUL.scala 102:19]
    .io_x1(m_1934_io_x1),
    .io_x2(m_1934_io_x2),
    .io_x3(m_1934_io_x3),
    .io_s(m_1934_io_s),
    .io_cout(m_1934_io_cout)
  );
  Adder m_1935 ( // @[MUL.scala 102:19]
    .io_x1(m_1935_io_x1),
    .io_x2(m_1935_io_x2),
    .io_x3(m_1935_io_x3),
    .io_s(m_1935_io_s),
    .io_cout(m_1935_io_cout)
  );
  Adder m_1936 ( // @[MUL.scala 102:19]
    .io_x1(m_1936_io_x1),
    .io_x2(m_1936_io_x2),
    .io_x3(m_1936_io_x3),
    .io_s(m_1936_io_s),
    .io_cout(m_1936_io_cout)
  );
  Adder m_1937 ( // @[MUL.scala 102:19]
    .io_x1(m_1937_io_x1),
    .io_x2(m_1937_io_x2),
    .io_x3(m_1937_io_x3),
    .io_s(m_1937_io_s),
    .io_cout(m_1937_io_cout)
  );
  Adder m_1938 ( // @[MUL.scala 102:19]
    .io_x1(m_1938_io_x1),
    .io_x2(m_1938_io_x2),
    .io_x3(m_1938_io_x3),
    .io_s(m_1938_io_s),
    .io_cout(m_1938_io_cout)
  );
  Adder m_1939 ( // @[MUL.scala 102:19]
    .io_x1(m_1939_io_x1),
    .io_x2(m_1939_io_x2),
    .io_x3(m_1939_io_x3),
    .io_s(m_1939_io_s),
    .io_cout(m_1939_io_cout)
  );
  Adder m_1940 ( // @[MUL.scala 102:19]
    .io_x1(m_1940_io_x1),
    .io_x2(m_1940_io_x2),
    .io_x3(m_1940_io_x3),
    .io_s(m_1940_io_s),
    .io_cout(m_1940_io_cout)
  );
  Adder m_1941 ( // @[MUL.scala 102:19]
    .io_x1(m_1941_io_x1),
    .io_x2(m_1941_io_x2),
    .io_x3(m_1941_io_x3),
    .io_s(m_1941_io_s),
    .io_cout(m_1941_io_cout)
  );
  Adder m_1942 ( // @[MUL.scala 102:19]
    .io_x1(m_1942_io_x1),
    .io_x2(m_1942_io_x2),
    .io_x3(m_1942_io_x3),
    .io_s(m_1942_io_s),
    .io_cout(m_1942_io_cout)
  );
  Adder m_1943 ( // @[MUL.scala 102:19]
    .io_x1(m_1943_io_x1),
    .io_x2(m_1943_io_x2),
    .io_x3(m_1943_io_x3),
    .io_s(m_1943_io_s),
    .io_cout(m_1943_io_cout)
  );
  Half_Adder m_1944 ( // @[MUL.scala 124:19]
    .io_in_0(m_1944_io_in_0),
    .io_in_1(m_1944_io_in_1),
    .io_out_0(m_1944_io_out_0),
    .io_out_1(m_1944_io_out_1)
  );
  Half_Adder m_1945 ( // @[MUL.scala 124:19]
    .io_in_0(m_1945_io_in_0),
    .io_in_1(m_1945_io_in_1),
    .io_out_0(m_1945_io_out_0),
    .io_out_1(m_1945_io_out_1)
  );
  Half_Adder m_1946 ( // @[MUL.scala 124:19]
    .io_in_0(m_1946_io_in_0),
    .io_in_1(m_1946_io_in_1),
    .io_out_0(m_1946_io_out_0),
    .io_out_1(m_1946_io_out_1)
  );
  Half_Adder m_1947 ( // @[MUL.scala 124:19]
    .io_in_0(m_1947_io_in_0),
    .io_in_1(m_1947_io_in_1),
    .io_out_0(m_1947_io_out_0),
    .io_out_1(m_1947_io_out_1)
  );
  Half_Adder m_1948 ( // @[MUL.scala 124:19]
    .io_in_0(m_1948_io_in_0),
    .io_in_1(m_1948_io_in_1),
    .io_out_0(m_1948_io_out_0),
    .io_out_1(m_1948_io_out_1)
  );
  Half_Adder m_1949 ( // @[MUL.scala 124:19]
    .io_in_0(m_1949_io_in_0),
    .io_in_1(m_1949_io_in_1),
    .io_out_0(m_1949_io_out_0),
    .io_out_1(m_1949_io_out_1)
  );
  Half_Adder m_1950 ( // @[MUL.scala 124:19]
    .io_in_0(m_1950_io_in_0),
    .io_in_1(m_1950_io_in_1),
    .io_out_0(m_1950_io_out_0),
    .io_out_1(m_1950_io_out_1)
  );
  Half_Adder m_1951 ( // @[MUL.scala 124:19]
    .io_in_0(m_1951_io_in_0),
    .io_in_1(m_1951_io_in_1),
    .io_out_0(m_1951_io_out_0),
    .io_out_1(m_1951_io_out_1)
  );
  Half_Adder m_1952 ( // @[MUL.scala 124:19]
    .io_in_0(m_1952_io_in_0),
    .io_in_1(m_1952_io_in_1),
    .io_out_0(m_1952_io_out_0),
    .io_out_1(m_1952_io_out_1)
  );
  Half_Adder m_1953 ( // @[MUL.scala 124:19]
    .io_in_0(m_1953_io_in_0),
    .io_in_1(m_1953_io_in_1),
    .io_out_0(m_1953_io_out_0),
    .io_out_1(m_1953_io_out_1)
  );
  Half_Adder m_1954 ( // @[MUL.scala 124:19]
    .io_in_0(m_1954_io_in_0),
    .io_in_1(m_1954_io_in_1),
    .io_out_0(m_1954_io_out_0),
    .io_out_1(m_1954_io_out_1)
  );
  Half_Adder m_1955 ( // @[MUL.scala 124:19]
    .io_in_0(m_1955_io_in_0),
    .io_in_1(m_1955_io_in_1),
    .io_out_0(m_1955_io_out_0),
    .io_out_1(m_1955_io_out_1)
  );
  Half_Adder m_1956 ( // @[MUL.scala 124:19]
    .io_in_0(m_1956_io_in_0),
    .io_in_1(m_1956_io_in_1),
    .io_out_0(m_1956_io_out_0),
    .io_out_1(m_1956_io_out_1)
  );
  Half_Adder m_1957 ( // @[MUL.scala 124:19]
    .io_in_0(m_1957_io_in_0),
    .io_in_1(m_1957_io_in_1),
    .io_out_0(m_1957_io_out_0),
    .io_out_1(m_1957_io_out_1)
  );
  Half_Adder m_1958 ( // @[MUL.scala 124:19]
    .io_in_0(m_1958_io_in_0),
    .io_in_1(m_1958_io_in_1),
    .io_out_0(m_1958_io_out_0),
    .io_out_1(m_1958_io_out_1)
  );
  Half_Adder m_1959 ( // @[MUL.scala 124:19]
    .io_in_0(m_1959_io_in_0),
    .io_in_1(m_1959_io_in_1),
    .io_out_0(m_1959_io_out_0),
    .io_out_1(m_1959_io_out_1)
  );
  Half_Adder m_1960 ( // @[MUL.scala 124:19]
    .io_in_0(m_1960_io_in_0),
    .io_in_1(m_1960_io_in_1),
    .io_out_0(m_1960_io_out_0),
    .io_out_1(m_1960_io_out_1)
  );
  Half_Adder m_1961 ( // @[MUL.scala 124:19]
    .io_in_0(m_1961_io_in_0),
    .io_in_1(m_1961_io_in_1),
    .io_out_0(m_1961_io_out_0),
    .io_out_1(m_1961_io_out_1)
  );
  Half_Adder m_1962 ( // @[MUL.scala 124:19]
    .io_in_0(m_1962_io_in_0),
    .io_in_1(m_1962_io_in_1),
    .io_out_0(m_1962_io_out_0),
    .io_out_1(m_1962_io_out_1)
  );
  Half_Adder m_1963 ( // @[MUL.scala 124:19]
    .io_in_0(m_1963_io_in_0),
    .io_in_1(m_1963_io_in_1),
    .io_out_0(m_1963_io_out_0),
    .io_out_1(m_1963_io_out_1)
  );
  Half_Adder m_1964 ( // @[MUL.scala 124:19]
    .io_in_0(m_1964_io_in_0),
    .io_in_1(m_1964_io_in_1),
    .io_out_0(m_1964_io_out_0),
    .io_out_1(m_1964_io_out_1)
  );
  Half_Adder m_1965 ( // @[MUL.scala 124:19]
    .io_in_0(m_1965_io_in_0),
    .io_in_1(m_1965_io_in_1),
    .io_out_0(m_1965_io_out_0),
    .io_out_1(m_1965_io_out_1)
  );
  Half_Adder m_1966 ( // @[MUL.scala 124:19]
    .io_in_0(m_1966_io_in_0),
    .io_in_1(m_1966_io_in_1),
    .io_out_0(m_1966_io_out_0),
    .io_out_1(m_1966_io_out_1)
  );
  Adder m_1967 ( // @[MUL.scala 102:19]
    .io_x1(m_1967_io_x1),
    .io_x2(m_1967_io_x2),
    .io_x3(m_1967_io_x3),
    .io_s(m_1967_io_s),
    .io_cout(m_1967_io_cout)
  );
  Adder m_1968 ( // @[MUL.scala 102:19]
    .io_x1(m_1968_io_x1),
    .io_x2(m_1968_io_x2),
    .io_x3(m_1968_io_x3),
    .io_s(m_1968_io_s),
    .io_cout(m_1968_io_cout)
  );
  Adder m_1969 ( // @[MUL.scala 102:19]
    .io_x1(m_1969_io_x1),
    .io_x2(m_1969_io_x2),
    .io_x3(m_1969_io_x3),
    .io_s(m_1969_io_s),
    .io_cout(m_1969_io_cout)
  );
  Adder m_1970 ( // @[MUL.scala 102:19]
    .io_x1(m_1970_io_x1),
    .io_x2(m_1970_io_x2),
    .io_x3(m_1970_io_x3),
    .io_s(m_1970_io_s),
    .io_cout(m_1970_io_cout)
  );
  Adder m_1971 ( // @[MUL.scala 102:19]
    .io_x1(m_1971_io_x1),
    .io_x2(m_1971_io_x2),
    .io_x3(m_1971_io_x3),
    .io_s(m_1971_io_s),
    .io_cout(m_1971_io_cout)
  );
  Adder m_1972 ( // @[MUL.scala 102:19]
    .io_x1(m_1972_io_x1),
    .io_x2(m_1972_io_x2),
    .io_x3(m_1972_io_x3),
    .io_s(m_1972_io_s),
    .io_cout(m_1972_io_cout)
  );
  Adder m_1973 ( // @[MUL.scala 102:19]
    .io_x1(m_1973_io_x1),
    .io_x2(m_1973_io_x2),
    .io_x3(m_1973_io_x3),
    .io_s(m_1973_io_s),
    .io_cout(m_1973_io_cout)
  );
  Adder m_1974 ( // @[MUL.scala 102:19]
    .io_x1(m_1974_io_x1),
    .io_x2(m_1974_io_x2),
    .io_x3(m_1974_io_x3),
    .io_s(m_1974_io_s),
    .io_cout(m_1974_io_cout)
  );
  Adder m_1975 ( // @[MUL.scala 102:19]
    .io_x1(m_1975_io_x1),
    .io_x2(m_1975_io_x2),
    .io_x3(m_1975_io_x3),
    .io_s(m_1975_io_s),
    .io_cout(m_1975_io_cout)
  );
  Adder m_1976 ( // @[MUL.scala 102:19]
    .io_x1(m_1976_io_x1),
    .io_x2(m_1976_io_x2),
    .io_x3(m_1976_io_x3),
    .io_s(m_1976_io_s),
    .io_cout(m_1976_io_cout)
  );
  Adder m_1977 ( // @[MUL.scala 102:19]
    .io_x1(m_1977_io_x1),
    .io_x2(m_1977_io_x2),
    .io_x3(m_1977_io_x3),
    .io_s(m_1977_io_s),
    .io_cout(m_1977_io_cout)
  );
  Adder m_1978 ( // @[MUL.scala 102:19]
    .io_x1(m_1978_io_x1),
    .io_x2(m_1978_io_x2),
    .io_x3(m_1978_io_x3),
    .io_s(m_1978_io_s),
    .io_cout(m_1978_io_cout)
  );
  Adder m_1979 ( // @[MUL.scala 102:19]
    .io_x1(m_1979_io_x1),
    .io_x2(m_1979_io_x2),
    .io_x3(m_1979_io_x3),
    .io_s(m_1979_io_s),
    .io_cout(m_1979_io_cout)
  );
  Adder m_1980 ( // @[MUL.scala 102:19]
    .io_x1(m_1980_io_x1),
    .io_x2(m_1980_io_x2),
    .io_x3(m_1980_io_x3),
    .io_s(m_1980_io_s),
    .io_cout(m_1980_io_cout)
  );
  Adder m_1981 ( // @[MUL.scala 102:19]
    .io_x1(m_1981_io_x1),
    .io_x2(m_1981_io_x2),
    .io_x3(m_1981_io_x3),
    .io_s(m_1981_io_s),
    .io_cout(m_1981_io_cout)
  );
  Adder m_1982 ( // @[MUL.scala 102:19]
    .io_x1(m_1982_io_x1),
    .io_x2(m_1982_io_x2),
    .io_x3(m_1982_io_x3),
    .io_s(m_1982_io_s),
    .io_cout(m_1982_io_cout)
  );
  Adder m_1983 ( // @[MUL.scala 102:19]
    .io_x1(m_1983_io_x1),
    .io_x2(m_1983_io_x2),
    .io_x3(m_1983_io_x3),
    .io_s(m_1983_io_s),
    .io_cout(m_1983_io_cout)
  );
  Adder m_1984 ( // @[MUL.scala 102:19]
    .io_x1(m_1984_io_x1),
    .io_x2(m_1984_io_x2),
    .io_x3(m_1984_io_x3),
    .io_s(m_1984_io_s),
    .io_cout(m_1984_io_cout)
  );
  Adder m_1985 ( // @[MUL.scala 102:19]
    .io_x1(m_1985_io_x1),
    .io_x2(m_1985_io_x2),
    .io_x3(m_1985_io_x3),
    .io_s(m_1985_io_s),
    .io_cout(m_1985_io_cout)
  );
  Adder m_1986 ( // @[MUL.scala 102:19]
    .io_x1(m_1986_io_x1),
    .io_x2(m_1986_io_x2),
    .io_x3(m_1986_io_x3),
    .io_s(m_1986_io_s),
    .io_cout(m_1986_io_cout)
  );
  Adder m_1987 ( // @[MUL.scala 102:19]
    .io_x1(m_1987_io_x1),
    .io_x2(m_1987_io_x2),
    .io_x3(m_1987_io_x3),
    .io_s(m_1987_io_s),
    .io_cout(m_1987_io_cout)
  );
  Adder m_1988 ( // @[MUL.scala 102:19]
    .io_x1(m_1988_io_x1),
    .io_x2(m_1988_io_x2),
    .io_x3(m_1988_io_x3),
    .io_s(m_1988_io_s),
    .io_cout(m_1988_io_cout)
  );
  Half_Adder m_1989 ( // @[MUL.scala 124:19]
    .io_in_0(m_1989_io_in_0),
    .io_in_1(m_1989_io_in_1),
    .io_out_0(m_1989_io_out_0),
    .io_out_1(m_1989_io_out_1)
  );
  Adder m_1990 ( // @[MUL.scala 102:19]
    .io_x1(m_1990_io_x1),
    .io_x2(m_1990_io_x2),
    .io_x3(m_1990_io_x3),
    .io_s(m_1990_io_s),
    .io_cout(m_1990_io_cout)
  );
  Half_Adder m_1991 ( // @[MUL.scala 124:19]
    .io_in_0(m_1991_io_in_0),
    .io_in_1(m_1991_io_in_1),
    .io_out_0(m_1991_io_out_0),
    .io_out_1(m_1991_io_out_1)
  );
  Adder m_1992 ( // @[MUL.scala 102:19]
    .io_x1(m_1992_io_x1),
    .io_x2(m_1992_io_x2),
    .io_x3(m_1992_io_x3),
    .io_s(m_1992_io_s),
    .io_cout(m_1992_io_cout)
  );
  Half_Adder m_1993 ( // @[MUL.scala 124:19]
    .io_in_0(m_1993_io_in_0),
    .io_in_1(m_1993_io_in_1),
    .io_out_0(m_1993_io_out_0),
    .io_out_1(m_1993_io_out_1)
  );
  Adder m_1994 ( // @[MUL.scala 102:19]
    .io_x1(m_1994_io_x1),
    .io_x2(m_1994_io_x2),
    .io_x3(m_1994_io_x3),
    .io_s(m_1994_io_s),
    .io_cout(m_1994_io_cout)
  );
  Half_Adder m_1995 ( // @[MUL.scala 124:19]
    .io_in_0(m_1995_io_in_0),
    .io_in_1(m_1995_io_in_1),
    .io_out_0(m_1995_io_out_0),
    .io_out_1(m_1995_io_out_1)
  );
  Adder m_1996 ( // @[MUL.scala 102:19]
    .io_x1(m_1996_io_x1),
    .io_x2(m_1996_io_x2),
    .io_x3(m_1996_io_x3),
    .io_s(m_1996_io_s),
    .io_cout(m_1996_io_cout)
  );
  Half_Adder m_1997 ( // @[MUL.scala 124:19]
    .io_in_0(m_1997_io_in_0),
    .io_in_1(m_1997_io_in_1),
    .io_out_0(m_1997_io_out_0),
    .io_out_1(m_1997_io_out_1)
  );
  Adder m_1998 ( // @[MUL.scala 102:19]
    .io_x1(m_1998_io_x1),
    .io_x2(m_1998_io_x2),
    .io_x3(m_1998_io_x3),
    .io_s(m_1998_io_s),
    .io_cout(m_1998_io_cout)
  );
  Half_Adder m_1999 ( // @[MUL.scala 124:19]
    .io_in_0(m_1999_io_in_0),
    .io_in_1(m_1999_io_in_1),
    .io_out_0(m_1999_io_out_0),
    .io_out_1(m_1999_io_out_1)
  );
  Adder m_2000 ( // @[MUL.scala 102:19]
    .io_x1(m_2000_io_x1),
    .io_x2(m_2000_io_x2),
    .io_x3(m_2000_io_x3),
    .io_s(m_2000_io_s),
    .io_cout(m_2000_io_cout)
  );
  Half_Adder m_2001 ( // @[MUL.scala 124:19]
    .io_in_0(m_2001_io_in_0),
    .io_in_1(m_2001_io_in_1),
    .io_out_0(m_2001_io_out_0),
    .io_out_1(m_2001_io_out_1)
  );
  Adder m_2002 ( // @[MUL.scala 102:19]
    .io_x1(m_2002_io_x1),
    .io_x2(m_2002_io_x2),
    .io_x3(m_2002_io_x3),
    .io_s(m_2002_io_s),
    .io_cout(m_2002_io_cout)
  );
  Adder m_2003 ( // @[MUL.scala 102:19]
    .io_x1(m_2003_io_x1),
    .io_x2(m_2003_io_x2),
    .io_x3(m_2003_io_x3),
    .io_s(m_2003_io_s),
    .io_cout(m_2003_io_cout)
  );
  Adder m_2004 ( // @[MUL.scala 102:19]
    .io_x1(m_2004_io_x1),
    .io_x2(m_2004_io_x2),
    .io_x3(m_2004_io_x3),
    .io_s(m_2004_io_s),
    .io_cout(m_2004_io_cout)
  );
  Adder m_2005 ( // @[MUL.scala 102:19]
    .io_x1(m_2005_io_x1),
    .io_x2(m_2005_io_x2),
    .io_x3(m_2005_io_x3),
    .io_s(m_2005_io_s),
    .io_cout(m_2005_io_cout)
  );
  Adder m_2006 ( // @[MUL.scala 102:19]
    .io_x1(m_2006_io_x1),
    .io_x2(m_2006_io_x2),
    .io_x3(m_2006_io_x3),
    .io_s(m_2006_io_s),
    .io_cout(m_2006_io_cout)
  );
  Adder m_2007 ( // @[MUL.scala 102:19]
    .io_x1(m_2007_io_x1),
    .io_x2(m_2007_io_x2),
    .io_x3(m_2007_io_x3),
    .io_s(m_2007_io_s),
    .io_cout(m_2007_io_cout)
  );
  Adder m_2008 ( // @[MUL.scala 102:19]
    .io_x1(m_2008_io_x1),
    .io_x2(m_2008_io_x2),
    .io_x3(m_2008_io_x3),
    .io_s(m_2008_io_s),
    .io_cout(m_2008_io_cout)
  );
  Adder m_2009 ( // @[MUL.scala 102:19]
    .io_x1(m_2009_io_x1),
    .io_x2(m_2009_io_x2),
    .io_x3(m_2009_io_x3),
    .io_s(m_2009_io_s),
    .io_cout(m_2009_io_cout)
  );
  Adder m_2010 ( // @[MUL.scala 102:19]
    .io_x1(m_2010_io_x1),
    .io_x2(m_2010_io_x2),
    .io_x3(m_2010_io_x3),
    .io_s(m_2010_io_s),
    .io_cout(m_2010_io_cout)
  );
  Adder m_2011 ( // @[MUL.scala 102:19]
    .io_x1(m_2011_io_x1),
    .io_x2(m_2011_io_x2),
    .io_x3(m_2011_io_x3),
    .io_s(m_2011_io_s),
    .io_cout(m_2011_io_cout)
  );
  Adder m_2012 ( // @[MUL.scala 102:19]
    .io_x1(m_2012_io_x1),
    .io_x2(m_2012_io_x2),
    .io_x3(m_2012_io_x3),
    .io_s(m_2012_io_s),
    .io_cout(m_2012_io_cout)
  );
  Adder m_2013 ( // @[MUL.scala 102:19]
    .io_x1(m_2013_io_x1),
    .io_x2(m_2013_io_x2),
    .io_x3(m_2013_io_x3),
    .io_s(m_2013_io_s),
    .io_cout(m_2013_io_cout)
  );
  Adder m_2014 ( // @[MUL.scala 102:19]
    .io_x1(m_2014_io_x1),
    .io_x2(m_2014_io_x2),
    .io_x3(m_2014_io_x3),
    .io_s(m_2014_io_s),
    .io_cout(m_2014_io_cout)
  );
  Adder m_2015 ( // @[MUL.scala 102:19]
    .io_x1(m_2015_io_x1),
    .io_x2(m_2015_io_x2),
    .io_x3(m_2015_io_x3),
    .io_s(m_2015_io_s),
    .io_cout(m_2015_io_cout)
  );
  Adder m_2016 ( // @[MUL.scala 102:19]
    .io_x1(m_2016_io_x1),
    .io_x2(m_2016_io_x2),
    .io_x3(m_2016_io_x3),
    .io_s(m_2016_io_s),
    .io_cout(m_2016_io_cout)
  );
  Adder m_2017 ( // @[MUL.scala 102:19]
    .io_x1(m_2017_io_x1),
    .io_x2(m_2017_io_x2),
    .io_x3(m_2017_io_x3),
    .io_s(m_2017_io_s),
    .io_cout(m_2017_io_cout)
  );
  Adder m_2018 ( // @[MUL.scala 102:19]
    .io_x1(m_2018_io_x1),
    .io_x2(m_2018_io_x2),
    .io_x3(m_2018_io_x3),
    .io_s(m_2018_io_s),
    .io_cout(m_2018_io_cout)
  );
  Adder m_2019 ( // @[MUL.scala 102:19]
    .io_x1(m_2019_io_x1),
    .io_x2(m_2019_io_x2),
    .io_x3(m_2019_io_x3),
    .io_s(m_2019_io_s),
    .io_cout(m_2019_io_cout)
  );
  Adder m_2020 ( // @[MUL.scala 102:19]
    .io_x1(m_2020_io_x1),
    .io_x2(m_2020_io_x2),
    .io_x3(m_2020_io_x3),
    .io_s(m_2020_io_s),
    .io_cout(m_2020_io_cout)
  );
  Adder m_2021 ( // @[MUL.scala 102:19]
    .io_x1(m_2021_io_x1),
    .io_x2(m_2021_io_x2),
    .io_x3(m_2021_io_x3),
    .io_s(m_2021_io_s),
    .io_cout(m_2021_io_cout)
  );
  Adder m_2022 ( // @[MUL.scala 102:19]
    .io_x1(m_2022_io_x1),
    .io_x2(m_2022_io_x2),
    .io_x3(m_2022_io_x3),
    .io_s(m_2022_io_s),
    .io_cout(m_2022_io_cout)
  );
  Adder m_2023 ( // @[MUL.scala 102:19]
    .io_x1(m_2023_io_x1),
    .io_x2(m_2023_io_x2),
    .io_x3(m_2023_io_x3),
    .io_s(m_2023_io_s),
    .io_cout(m_2023_io_cout)
  );
  Adder m_2024 ( // @[MUL.scala 102:19]
    .io_x1(m_2024_io_x1),
    .io_x2(m_2024_io_x2),
    .io_x3(m_2024_io_x3),
    .io_s(m_2024_io_s),
    .io_cout(m_2024_io_cout)
  );
  Adder m_2025 ( // @[MUL.scala 102:19]
    .io_x1(m_2025_io_x1),
    .io_x2(m_2025_io_x2),
    .io_x3(m_2025_io_x3),
    .io_s(m_2025_io_s),
    .io_cout(m_2025_io_cout)
  );
  Adder m_2026 ( // @[MUL.scala 102:19]
    .io_x1(m_2026_io_x1),
    .io_x2(m_2026_io_x2),
    .io_x3(m_2026_io_x3),
    .io_s(m_2026_io_s),
    .io_cout(m_2026_io_cout)
  );
  Adder m_2027 ( // @[MUL.scala 102:19]
    .io_x1(m_2027_io_x1),
    .io_x2(m_2027_io_x2),
    .io_x3(m_2027_io_x3),
    .io_s(m_2027_io_s),
    .io_cout(m_2027_io_cout)
  );
  Adder m_2028 ( // @[MUL.scala 102:19]
    .io_x1(m_2028_io_x1),
    .io_x2(m_2028_io_x2),
    .io_x3(m_2028_io_x3),
    .io_s(m_2028_io_s),
    .io_cout(m_2028_io_cout)
  );
  Adder m_2029 ( // @[MUL.scala 102:19]
    .io_x1(m_2029_io_x1),
    .io_x2(m_2029_io_x2),
    .io_x3(m_2029_io_x3),
    .io_s(m_2029_io_s),
    .io_cout(m_2029_io_cout)
  );
  Adder m_2030 ( // @[MUL.scala 102:19]
    .io_x1(m_2030_io_x1),
    .io_x2(m_2030_io_x2),
    .io_x3(m_2030_io_x3),
    .io_s(m_2030_io_s),
    .io_cout(m_2030_io_cout)
  );
  Adder m_2031 ( // @[MUL.scala 102:19]
    .io_x1(m_2031_io_x1),
    .io_x2(m_2031_io_x2),
    .io_x3(m_2031_io_x3),
    .io_s(m_2031_io_s),
    .io_cout(m_2031_io_cout)
  );
  Adder m_2032 ( // @[MUL.scala 102:19]
    .io_x1(m_2032_io_x1),
    .io_x2(m_2032_io_x2),
    .io_x3(m_2032_io_x3),
    .io_s(m_2032_io_s),
    .io_cout(m_2032_io_cout)
  );
  Adder m_2033 ( // @[MUL.scala 102:19]
    .io_x1(m_2033_io_x1),
    .io_x2(m_2033_io_x2),
    .io_x3(m_2033_io_x3),
    .io_s(m_2033_io_s),
    .io_cout(m_2033_io_cout)
  );
  Adder m_2034 ( // @[MUL.scala 102:19]
    .io_x1(m_2034_io_x1),
    .io_x2(m_2034_io_x2),
    .io_x3(m_2034_io_x3),
    .io_s(m_2034_io_s),
    .io_cout(m_2034_io_cout)
  );
  Adder m_2035 ( // @[MUL.scala 102:19]
    .io_x1(m_2035_io_x1),
    .io_x2(m_2035_io_x2),
    .io_x3(m_2035_io_x3),
    .io_s(m_2035_io_s),
    .io_cout(m_2035_io_cout)
  );
  Adder m_2036 ( // @[MUL.scala 102:19]
    .io_x1(m_2036_io_x1),
    .io_x2(m_2036_io_x2),
    .io_x3(m_2036_io_x3),
    .io_s(m_2036_io_s),
    .io_cout(m_2036_io_cout)
  );
  Adder m_2037 ( // @[MUL.scala 102:19]
    .io_x1(m_2037_io_x1),
    .io_x2(m_2037_io_x2),
    .io_x3(m_2037_io_x3),
    .io_s(m_2037_io_s),
    .io_cout(m_2037_io_cout)
  );
  Adder m_2038 ( // @[MUL.scala 102:19]
    .io_x1(m_2038_io_x1),
    .io_x2(m_2038_io_x2),
    .io_x3(m_2038_io_x3),
    .io_s(m_2038_io_s),
    .io_cout(m_2038_io_cout)
  );
  Adder m_2039 ( // @[MUL.scala 102:19]
    .io_x1(m_2039_io_x1),
    .io_x2(m_2039_io_x2),
    .io_x3(m_2039_io_x3),
    .io_s(m_2039_io_s),
    .io_cout(m_2039_io_cout)
  );
  Adder m_2040 ( // @[MUL.scala 102:19]
    .io_x1(m_2040_io_x1),
    .io_x2(m_2040_io_x2),
    .io_x3(m_2040_io_x3),
    .io_s(m_2040_io_s),
    .io_cout(m_2040_io_cout)
  );
  Adder m_2041 ( // @[MUL.scala 102:19]
    .io_x1(m_2041_io_x1),
    .io_x2(m_2041_io_x2),
    .io_x3(m_2041_io_x3),
    .io_s(m_2041_io_s),
    .io_cout(m_2041_io_cout)
  );
  Adder m_2042 ( // @[MUL.scala 102:19]
    .io_x1(m_2042_io_x1),
    .io_x2(m_2042_io_x2),
    .io_x3(m_2042_io_x3),
    .io_s(m_2042_io_s),
    .io_cout(m_2042_io_cout)
  );
  Adder m_2043 ( // @[MUL.scala 102:19]
    .io_x1(m_2043_io_x1),
    .io_x2(m_2043_io_x2),
    .io_x3(m_2043_io_x3),
    .io_s(m_2043_io_s),
    .io_cout(m_2043_io_cout)
  );
  Adder m_2044 ( // @[MUL.scala 102:19]
    .io_x1(m_2044_io_x1),
    .io_x2(m_2044_io_x2),
    .io_x3(m_2044_io_x3),
    .io_s(m_2044_io_s),
    .io_cout(m_2044_io_cout)
  );
  Adder m_2045 ( // @[MUL.scala 102:19]
    .io_x1(m_2045_io_x1),
    .io_x2(m_2045_io_x2),
    .io_x3(m_2045_io_x3),
    .io_s(m_2045_io_s),
    .io_cout(m_2045_io_cout)
  );
  Adder m_2046 ( // @[MUL.scala 102:19]
    .io_x1(m_2046_io_x1),
    .io_x2(m_2046_io_x2),
    .io_x3(m_2046_io_x3),
    .io_s(m_2046_io_s),
    .io_cout(m_2046_io_cout)
  );
  Adder m_2047 ( // @[MUL.scala 102:19]
    .io_x1(m_2047_io_x1),
    .io_x2(m_2047_io_x2),
    .io_x3(m_2047_io_x3),
    .io_s(m_2047_io_s),
    .io_cout(m_2047_io_cout)
  );
  Adder m_2048 ( // @[MUL.scala 102:19]
    .io_x1(m_2048_io_x1),
    .io_x2(m_2048_io_x2),
    .io_x3(m_2048_io_x3),
    .io_s(m_2048_io_s),
    .io_cout(m_2048_io_cout)
  );
  Adder m_2049 ( // @[MUL.scala 102:19]
    .io_x1(m_2049_io_x1),
    .io_x2(m_2049_io_x2),
    .io_x3(m_2049_io_x3),
    .io_s(m_2049_io_s),
    .io_cout(m_2049_io_cout)
  );
  Adder m_2050 ( // @[MUL.scala 102:19]
    .io_x1(m_2050_io_x1),
    .io_x2(m_2050_io_x2),
    .io_x3(m_2050_io_x3),
    .io_s(m_2050_io_s),
    .io_cout(m_2050_io_cout)
  );
  Adder m_2051 ( // @[MUL.scala 102:19]
    .io_x1(m_2051_io_x1),
    .io_x2(m_2051_io_x2),
    .io_x3(m_2051_io_x3),
    .io_s(m_2051_io_s),
    .io_cout(m_2051_io_cout)
  );
  Adder m_2052 ( // @[MUL.scala 102:19]
    .io_x1(m_2052_io_x1),
    .io_x2(m_2052_io_x2),
    .io_x3(m_2052_io_x3),
    .io_s(m_2052_io_s),
    .io_cout(m_2052_io_cout)
  );
  Adder m_2053 ( // @[MUL.scala 102:19]
    .io_x1(m_2053_io_x1),
    .io_x2(m_2053_io_x2),
    .io_x3(m_2053_io_x3),
    .io_s(m_2053_io_s),
    .io_cout(m_2053_io_cout)
  );
  Adder m_2054 ( // @[MUL.scala 102:19]
    .io_x1(m_2054_io_x1),
    .io_x2(m_2054_io_x2),
    .io_x3(m_2054_io_x3),
    .io_s(m_2054_io_s),
    .io_cout(m_2054_io_cout)
  );
  Adder m_2055 ( // @[MUL.scala 102:19]
    .io_x1(m_2055_io_x1),
    .io_x2(m_2055_io_x2),
    .io_x3(m_2055_io_x3),
    .io_s(m_2055_io_s),
    .io_cout(m_2055_io_cout)
  );
  Adder m_2056 ( // @[MUL.scala 102:19]
    .io_x1(m_2056_io_x1),
    .io_x2(m_2056_io_x2),
    .io_x3(m_2056_io_x3),
    .io_s(m_2056_io_s),
    .io_cout(m_2056_io_cout)
  );
  Adder m_2057 ( // @[MUL.scala 102:19]
    .io_x1(m_2057_io_x1),
    .io_x2(m_2057_io_x2),
    .io_x3(m_2057_io_x3),
    .io_s(m_2057_io_s),
    .io_cout(m_2057_io_cout)
  );
  Adder m_2058 ( // @[MUL.scala 102:19]
    .io_x1(m_2058_io_x1),
    .io_x2(m_2058_io_x2),
    .io_x3(m_2058_io_x3),
    .io_s(m_2058_io_s),
    .io_cout(m_2058_io_cout)
  );
  Adder m_2059 ( // @[MUL.scala 102:19]
    .io_x1(m_2059_io_x1),
    .io_x2(m_2059_io_x2),
    .io_x3(m_2059_io_x3),
    .io_s(m_2059_io_s),
    .io_cout(m_2059_io_cout)
  );
  Adder m_2060 ( // @[MUL.scala 102:19]
    .io_x1(m_2060_io_x1),
    .io_x2(m_2060_io_x2),
    .io_x3(m_2060_io_x3),
    .io_s(m_2060_io_s),
    .io_cout(m_2060_io_cout)
  );
  Adder m_2061 ( // @[MUL.scala 102:19]
    .io_x1(m_2061_io_x1),
    .io_x2(m_2061_io_x2),
    .io_x3(m_2061_io_x3),
    .io_s(m_2061_io_s),
    .io_cout(m_2061_io_cout)
  );
  Adder m_2062 ( // @[MUL.scala 102:19]
    .io_x1(m_2062_io_x1),
    .io_x2(m_2062_io_x2),
    .io_x3(m_2062_io_x3),
    .io_s(m_2062_io_s),
    .io_cout(m_2062_io_cout)
  );
  Adder m_2063 ( // @[MUL.scala 102:19]
    .io_x1(m_2063_io_x1),
    .io_x2(m_2063_io_x2),
    .io_x3(m_2063_io_x3),
    .io_s(m_2063_io_s),
    .io_cout(m_2063_io_cout)
  );
  Adder m_2064 ( // @[MUL.scala 102:19]
    .io_x1(m_2064_io_x1),
    .io_x2(m_2064_io_x2),
    .io_x3(m_2064_io_x3),
    .io_s(m_2064_io_s),
    .io_cout(m_2064_io_cout)
  );
  Adder m_2065 ( // @[MUL.scala 102:19]
    .io_x1(m_2065_io_x1),
    .io_x2(m_2065_io_x2),
    .io_x3(m_2065_io_x3),
    .io_s(m_2065_io_s),
    .io_cout(m_2065_io_cout)
  );
  Adder m_2066 ( // @[MUL.scala 102:19]
    .io_x1(m_2066_io_x1),
    .io_x2(m_2066_io_x2),
    .io_x3(m_2066_io_x3),
    .io_s(m_2066_io_s),
    .io_cout(m_2066_io_cout)
  );
  Adder m_2067 ( // @[MUL.scala 102:19]
    .io_x1(m_2067_io_x1),
    .io_x2(m_2067_io_x2),
    .io_x3(m_2067_io_x3),
    .io_s(m_2067_io_s),
    .io_cout(m_2067_io_cout)
  );
  Adder m_2068 ( // @[MUL.scala 102:19]
    .io_x1(m_2068_io_x1),
    .io_x2(m_2068_io_x2),
    .io_x3(m_2068_io_x3),
    .io_s(m_2068_io_s),
    .io_cout(m_2068_io_cout)
  );
  Adder m_2069 ( // @[MUL.scala 102:19]
    .io_x1(m_2069_io_x1),
    .io_x2(m_2069_io_x2),
    .io_x3(m_2069_io_x3),
    .io_s(m_2069_io_s),
    .io_cout(m_2069_io_cout)
  );
  Adder m_2070 ( // @[MUL.scala 102:19]
    .io_x1(m_2070_io_x1),
    .io_x2(m_2070_io_x2),
    .io_x3(m_2070_io_x3),
    .io_s(m_2070_io_s),
    .io_cout(m_2070_io_cout)
  );
  Adder m_2071 ( // @[MUL.scala 102:19]
    .io_x1(m_2071_io_x1),
    .io_x2(m_2071_io_x2),
    .io_x3(m_2071_io_x3),
    .io_s(m_2071_io_s),
    .io_cout(m_2071_io_cout)
  );
  Adder m_2072 ( // @[MUL.scala 102:19]
    .io_x1(m_2072_io_x1),
    .io_x2(m_2072_io_x2),
    .io_x3(m_2072_io_x3),
    .io_s(m_2072_io_s),
    .io_cout(m_2072_io_cout)
  );
  Adder m_2073 ( // @[MUL.scala 102:19]
    .io_x1(m_2073_io_x1),
    .io_x2(m_2073_io_x2),
    .io_x3(m_2073_io_x3),
    .io_s(m_2073_io_s),
    .io_cout(m_2073_io_cout)
  );
  Adder m_2074 ( // @[MUL.scala 102:19]
    .io_x1(m_2074_io_x1),
    .io_x2(m_2074_io_x2),
    .io_x3(m_2074_io_x3),
    .io_s(m_2074_io_s),
    .io_cout(m_2074_io_cout)
  );
  Adder m_2075 ( // @[MUL.scala 102:19]
    .io_x1(m_2075_io_x1),
    .io_x2(m_2075_io_x2),
    .io_x3(m_2075_io_x3),
    .io_s(m_2075_io_s),
    .io_cout(m_2075_io_cout)
  );
  Adder m_2076 ( // @[MUL.scala 102:19]
    .io_x1(m_2076_io_x1),
    .io_x2(m_2076_io_x2),
    .io_x3(m_2076_io_x3),
    .io_s(m_2076_io_s),
    .io_cout(m_2076_io_cout)
  );
  Adder m_2077 ( // @[MUL.scala 102:19]
    .io_x1(m_2077_io_x1),
    .io_x2(m_2077_io_x2),
    .io_x3(m_2077_io_x3),
    .io_s(m_2077_io_s),
    .io_cout(m_2077_io_cout)
  );
  Adder m_2078 ( // @[MUL.scala 102:19]
    .io_x1(m_2078_io_x1),
    .io_x2(m_2078_io_x2),
    .io_x3(m_2078_io_x3),
    .io_s(m_2078_io_s),
    .io_cout(m_2078_io_cout)
  );
  Adder m_2079 ( // @[MUL.scala 102:19]
    .io_x1(m_2079_io_x1),
    .io_x2(m_2079_io_x2),
    .io_x3(m_2079_io_x3),
    .io_s(m_2079_io_s),
    .io_cout(m_2079_io_cout)
  );
  Adder m_2080 ( // @[MUL.scala 102:19]
    .io_x1(m_2080_io_x1),
    .io_x2(m_2080_io_x2),
    .io_x3(m_2080_io_x3),
    .io_s(m_2080_io_s),
    .io_cout(m_2080_io_cout)
  );
  Adder m_2081 ( // @[MUL.scala 102:19]
    .io_x1(m_2081_io_x1),
    .io_x2(m_2081_io_x2),
    .io_x3(m_2081_io_x3),
    .io_s(m_2081_io_s),
    .io_cout(m_2081_io_cout)
  );
  Adder m_2082 ( // @[MUL.scala 102:19]
    .io_x1(m_2082_io_x1),
    .io_x2(m_2082_io_x2),
    .io_x3(m_2082_io_x3),
    .io_s(m_2082_io_s),
    .io_cout(m_2082_io_cout)
  );
  Adder m_2083 ( // @[MUL.scala 102:19]
    .io_x1(m_2083_io_x1),
    .io_x2(m_2083_io_x2),
    .io_x3(m_2083_io_x3),
    .io_s(m_2083_io_s),
    .io_cout(m_2083_io_cout)
  );
  Adder m_2084 ( // @[MUL.scala 102:19]
    .io_x1(m_2084_io_x1),
    .io_x2(m_2084_io_x2),
    .io_x3(m_2084_io_x3),
    .io_s(m_2084_io_s),
    .io_cout(m_2084_io_cout)
  );
  Adder m_2085 ( // @[MUL.scala 102:19]
    .io_x1(m_2085_io_x1),
    .io_x2(m_2085_io_x2),
    .io_x3(m_2085_io_x3),
    .io_s(m_2085_io_s),
    .io_cout(m_2085_io_cout)
  );
  Adder m_2086 ( // @[MUL.scala 102:19]
    .io_x1(m_2086_io_x1),
    .io_x2(m_2086_io_x2),
    .io_x3(m_2086_io_x3),
    .io_s(m_2086_io_s),
    .io_cout(m_2086_io_cout)
  );
  Adder m_2087 ( // @[MUL.scala 102:19]
    .io_x1(m_2087_io_x1),
    .io_x2(m_2087_io_x2),
    .io_x3(m_2087_io_x3),
    .io_s(m_2087_io_s),
    .io_cout(m_2087_io_cout)
  );
  Adder m_2088 ( // @[MUL.scala 102:19]
    .io_x1(m_2088_io_x1),
    .io_x2(m_2088_io_x2),
    .io_x3(m_2088_io_x3),
    .io_s(m_2088_io_s),
    .io_cout(m_2088_io_cout)
  );
  Adder m_2089 ( // @[MUL.scala 102:19]
    .io_x1(m_2089_io_x1),
    .io_x2(m_2089_io_x2),
    .io_x3(m_2089_io_x3),
    .io_s(m_2089_io_s),
    .io_cout(m_2089_io_cout)
  );
  Adder m_2090 ( // @[MUL.scala 102:19]
    .io_x1(m_2090_io_x1),
    .io_x2(m_2090_io_x2),
    .io_x3(m_2090_io_x3),
    .io_s(m_2090_io_s),
    .io_cout(m_2090_io_cout)
  );
  Adder m_2091 ( // @[MUL.scala 102:19]
    .io_x1(m_2091_io_x1),
    .io_x2(m_2091_io_x2),
    .io_x3(m_2091_io_x3),
    .io_s(m_2091_io_s),
    .io_cout(m_2091_io_cout)
  );
  Adder m_2092 ( // @[MUL.scala 102:19]
    .io_x1(m_2092_io_x1),
    .io_x2(m_2092_io_x2),
    .io_x3(m_2092_io_x3),
    .io_s(m_2092_io_s),
    .io_cout(m_2092_io_cout)
  );
  Adder m_2093 ( // @[MUL.scala 102:19]
    .io_x1(m_2093_io_x1),
    .io_x2(m_2093_io_x2),
    .io_x3(m_2093_io_x3),
    .io_s(m_2093_io_s),
    .io_cout(m_2093_io_cout)
  );
  Adder m_2094 ( // @[MUL.scala 102:19]
    .io_x1(m_2094_io_x1),
    .io_x2(m_2094_io_x2),
    .io_x3(m_2094_io_x3),
    .io_s(m_2094_io_s),
    .io_cout(m_2094_io_cout)
  );
  Half_Adder m_2095 ( // @[MUL.scala 124:19]
    .io_in_0(m_2095_io_in_0),
    .io_in_1(m_2095_io_in_1),
    .io_out_0(m_2095_io_out_0),
    .io_out_1(m_2095_io_out_1)
  );
  Adder m_2096 ( // @[MUL.scala 102:19]
    .io_x1(m_2096_io_x1),
    .io_x2(m_2096_io_x2),
    .io_x3(m_2096_io_x3),
    .io_s(m_2096_io_s),
    .io_cout(m_2096_io_cout)
  );
  Half_Adder m_2097 ( // @[MUL.scala 124:19]
    .io_in_0(m_2097_io_in_0),
    .io_in_1(m_2097_io_in_1),
    .io_out_0(m_2097_io_out_0),
    .io_out_1(m_2097_io_out_1)
  );
  Adder m_2098 ( // @[MUL.scala 102:19]
    .io_x1(m_2098_io_x1),
    .io_x2(m_2098_io_x2),
    .io_x3(m_2098_io_x3),
    .io_s(m_2098_io_s),
    .io_cout(m_2098_io_cout)
  );
  Half_Adder m_2099 ( // @[MUL.scala 124:19]
    .io_in_0(m_2099_io_in_0),
    .io_in_1(m_2099_io_in_1),
    .io_out_0(m_2099_io_out_0),
    .io_out_1(m_2099_io_out_1)
  );
  Adder m_2100 ( // @[MUL.scala 102:19]
    .io_x1(m_2100_io_x1),
    .io_x2(m_2100_io_x2),
    .io_x3(m_2100_io_x3),
    .io_s(m_2100_io_s),
    .io_cout(m_2100_io_cout)
  );
  Half_Adder m_2101 ( // @[MUL.scala 124:19]
    .io_in_0(m_2101_io_in_0),
    .io_in_1(m_2101_io_in_1),
    .io_out_0(m_2101_io_out_0),
    .io_out_1(m_2101_io_out_1)
  );
  Adder m_2102 ( // @[MUL.scala 102:19]
    .io_x1(m_2102_io_x1),
    .io_x2(m_2102_io_x2),
    .io_x3(m_2102_io_x3),
    .io_s(m_2102_io_s),
    .io_cout(m_2102_io_cout)
  );
  Half_Adder m_2103 ( // @[MUL.scala 124:19]
    .io_in_0(m_2103_io_in_0),
    .io_in_1(m_2103_io_in_1),
    .io_out_0(m_2103_io_out_0),
    .io_out_1(m_2103_io_out_1)
  );
  Adder m_2104 ( // @[MUL.scala 102:19]
    .io_x1(m_2104_io_x1),
    .io_x2(m_2104_io_x2),
    .io_x3(m_2104_io_x3),
    .io_s(m_2104_io_s),
    .io_cout(m_2104_io_cout)
  );
  Adder m_2105 ( // @[MUL.scala 102:19]
    .io_x1(m_2105_io_x1),
    .io_x2(m_2105_io_x2),
    .io_x3(m_2105_io_x3),
    .io_s(m_2105_io_s),
    .io_cout(m_2105_io_cout)
  );
  Adder m_2106 ( // @[MUL.scala 102:19]
    .io_x1(m_2106_io_x1),
    .io_x2(m_2106_io_x2),
    .io_x3(m_2106_io_x3),
    .io_s(m_2106_io_s),
    .io_cout(m_2106_io_cout)
  );
  Adder m_2107 ( // @[MUL.scala 102:19]
    .io_x1(m_2107_io_x1),
    .io_x2(m_2107_io_x2),
    .io_x3(m_2107_io_x3),
    .io_s(m_2107_io_s),
    .io_cout(m_2107_io_cout)
  );
  Adder m_2108 ( // @[MUL.scala 102:19]
    .io_x1(m_2108_io_x1),
    .io_x2(m_2108_io_x2),
    .io_x3(m_2108_io_x3),
    .io_s(m_2108_io_s),
    .io_cout(m_2108_io_cout)
  );
  Adder m_2109 ( // @[MUL.scala 102:19]
    .io_x1(m_2109_io_x1),
    .io_x2(m_2109_io_x2),
    .io_x3(m_2109_io_x3),
    .io_s(m_2109_io_s),
    .io_cout(m_2109_io_cout)
  );
  Adder m_2110 ( // @[MUL.scala 102:19]
    .io_x1(m_2110_io_x1),
    .io_x2(m_2110_io_x2),
    .io_x3(m_2110_io_x3),
    .io_s(m_2110_io_s),
    .io_cout(m_2110_io_cout)
  );
  Adder m_2111 ( // @[MUL.scala 102:19]
    .io_x1(m_2111_io_x1),
    .io_x2(m_2111_io_x2),
    .io_x3(m_2111_io_x3),
    .io_s(m_2111_io_s),
    .io_cout(m_2111_io_cout)
  );
  Adder m_2112 ( // @[MUL.scala 102:19]
    .io_x1(m_2112_io_x1),
    .io_x2(m_2112_io_x2),
    .io_x3(m_2112_io_x3),
    .io_s(m_2112_io_s),
    .io_cout(m_2112_io_cout)
  );
  Adder m_2113 ( // @[MUL.scala 102:19]
    .io_x1(m_2113_io_x1),
    .io_x2(m_2113_io_x2),
    .io_x3(m_2113_io_x3),
    .io_s(m_2113_io_s),
    .io_cout(m_2113_io_cout)
  );
  Adder m_2114 ( // @[MUL.scala 102:19]
    .io_x1(m_2114_io_x1),
    .io_x2(m_2114_io_x2),
    .io_x3(m_2114_io_x3),
    .io_s(m_2114_io_s),
    .io_cout(m_2114_io_cout)
  );
  Adder m_2115 ( // @[MUL.scala 102:19]
    .io_x1(m_2115_io_x1),
    .io_x2(m_2115_io_x2),
    .io_x3(m_2115_io_x3),
    .io_s(m_2115_io_s),
    .io_cout(m_2115_io_cout)
  );
  Adder m_2116 ( // @[MUL.scala 102:19]
    .io_x1(m_2116_io_x1),
    .io_x2(m_2116_io_x2),
    .io_x3(m_2116_io_x3),
    .io_s(m_2116_io_s),
    .io_cout(m_2116_io_cout)
  );
  Adder m_2117 ( // @[MUL.scala 102:19]
    .io_x1(m_2117_io_x1),
    .io_x2(m_2117_io_x2),
    .io_x3(m_2117_io_x3),
    .io_s(m_2117_io_s),
    .io_cout(m_2117_io_cout)
  );
  Adder m_2118 ( // @[MUL.scala 102:19]
    .io_x1(m_2118_io_x1),
    .io_x2(m_2118_io_x2),
    .io_x3(m_2118_io_x3),
    .io_s(m_2118_io_s),
    .io_cout(m_2118_io_cout)
  );
  Adder m_2119 ( // @[MUL.scala 102:19]
    .io_x1(m_2119_io_x1),
    .io_x2(m_2119_io_x2),
    .io_x3(m_2119_io_x3),
    .io_s(m_2119_io_s),
    .io_cout(m_2119_io_cout)
  );
  Adder m_2120 ( // @[MUL.scala 102:19]
    .io_x1(m_2120_io_x1),
    .io_x2(m_2120_io_x2),
    .io_x3(m_2120_io_x3),
    .io_s(m_2120_io_s),
    .io_cout(m_2120_io_cout)
  );
  Adder m_2121 ( // @[MUL.scala 102:19]
    .io_x1(m_2121_io_x1),
    .io_x2(m_2121_io_x2),
    .io_x3(m_2121_io_x3),
    .io_s(m_2121_io_s),
    .io_cout(m_2121_io_cout)
  );
  Adder m_2122 ( // @[MUL.scala 102:19]
    .io_x1(m_2122_io_x1),
    .io_x2(m_2122_io_x2),
    .io_x3(m_2122_io_x3),
    .io_s(m_2122_io_s),
    .io_cout(m_2122_io_cout)
  );
  Half_Adder m_2123 ( // @[MUL.scala 124:19]
    .io_in_0(m_2123_io_in_0),
    .io_in_1(m_2123_io_in_1),
    .io_out_0(m_2123_io_out_0),
    .io_out_1(m_2123_io_out_1)
  );
  Half_Adder m_2124 ( // @[MUL.scala 124:19]
    .io_in_0(m_2124_io_in_0),
    .io_in_1(m_2124_io_in_1),
    .io_out_0(m_2124_io_out_0),
    .io_out_1(m_2124_io_out_1)
  );
  Half_Adder m_2125 ( // @[MUL.scala 124:19]
    .io_in_0(m_2125_io_in_0),
    .io_in_1(m_2125_io_in_1),
    .io_out_0(m_2125_io_out_0),
    .io_out_1(m_2125_io_out_1)
  );
  Half_Adder m_2126 ( // @[MUL.scala 124:19]
    .io_in_0(m_2126_io_in_0),
    .io_in_1(m_2126_io_in_1),
    .io_out_0(m_2126_io_out_0),
    .io_out_1(m_2126_io_out_1)
  );
  Half_Adder m_2127 ( // @[MUL.scala 124:19]
    .io_in_0(m_2127_io_in_0),
    .io_in_1(m_2127_io_in_1),
    .io_out_0(m_2127_io_out_0),
    .io_out_1(m_2127_io_out_1)
  );
  Half_Adder m_2128 ( // @[MUL.scala 124:19]
    .io_in_0(m_2128_io_in_0),
    .io_in_1(m_2128_io_in_1),
    .io_out_0(m_2128_io_out_0),
    .io_out_1(m_2128_io_out_1)
  );
  Half_Adder m_2129 ( // @[MUL.scala 124:19]
    .io_in_0(m_2129_io_in_0),
    .io_in_1(m_2129_io_in_1),
    .io_out_0(m_2129_io_out_0),
    .io_out_1(m_2129_io_out_1)
  );
  Half_Adder m_2130 ( // @[MUL.scala 124:19]
    .io_in_0(m_2130_io_in_0),
    .io_in_1(m_2130_io_in_1),
    .io_out_0(m_2130_io_out_0),
    .io_out_1(m_2130_io_out_1)
  );
  Half_Adder m_2131 ( // @[MUL.scala 124:19]
    .io_in_0(m_2131_io_in_0),
    .io_in_1(m_2131_io_in_1),
    .io_out_0(m_2131_io_out_0),
    .io_out_1(m_2131_io_out_1)
  );
  Half_Adder m_2132 ( // @[MUL.scala 124:19]
    .io_in_0(m_2132_io_in_0),
    .io_in_1(m_2132_io_in_1),
    .io_out_0(m_2132_io_out_0),
    .io_out_1(m_2132_io_out_1)
  );
  Half_Adder m_2133 ( // @[MUL.scala 124:19]
    .io_in_0(m_2133_io_in_0),
    .io_in_1(m_2133_io_in_1),
    .io_out_0(m_2133_io_out_0),
    .io_out_1(m_2133_io_out_1)
  );
  Half_Adder m_2134 ( // @[MUL.scala 124:19]
    .io_in_0(m_2134_io_in_0),
    .io_in_1(m_2134_io_in_1),
    .io_out_0(m_2134_io_out_0),
    .io_out_1(m_2134_io_out_1)
  );
  Half_Adder m_2135 ( // @[MUL.scala 124:19]
    .io_in_0(m_2135_io_in_0),
    .io_in_1(m_2135_io_in_1),
    .io_out_0(m_2135_io_out_0),
    .io_out_1(m_2135_io_out_1)
  );
  Half_Adder m_2136 ( // @[MUL.scala 124:19]
    .io_in_0(m_2136_io_in_0),
    .io_in_1(m_2136_io_in_1),
    .io_out_0(m_2136_io_out_0),
    .io_out_1(m_2136_io_out_1)
  );
  Half_Adder m_2137 ( // @[MUL.scala 124:19]
    .io_in_0(m_2137_io_in_0),
    .io_in_1(m_2137_io_in_1),
    .io_out_0(m_2137_io_out_0),
    .io_out_1(m_2137_io_out_1)
  );
  Half_Adder m_2138 ( // @[MUL.scala 124:19]
    .io_in_0(m_2138_io_in_0),
    .io_in_1(m_2138_io_in_1),
    .io_out_0(m_2138_io_out_0),
    .io_out_1(m_2138_io_out_1)
  );
  Half_Adder m_2139 ( // @[MUL.scala 124:19]
    .io_in_0(m_2139_io_in_0),
    .io_in_1(m_2139_io_in_1),
    .io_out_0(m_2139_io_out_0),
    .io_out_1(m_2139_io_out_1)
  );
  Half_Adder m_2140 ( // @[MUL.scala 124:19]
    .io_in_0(m_2140_io_in_0),
    .io_in_1(m_2140_io_in_1),
    .io_out_0(m_2140_io_out_0),
    .io_out_1(m_2140_io_out_1)
  );
  Half_Adder m_2141 ( // @[MUL.scala 124:19]
    .io_in_0(m_2141_io_in_0),
    .io_in_1(m_2141_io_in_1),
    .io_out_0(m_2141_io_out_0),
    .io_out_1(m_2141_io_out_1)
  );
  Half_Adder m_2142 ( // @[MUL.scala 124:19]
    .io_in_0(m_2142_io_in_0),
    .io_in_1(m_2142_io_in_1),
    .io_out_0(m_2142_io_out_0),
    .io_out_1(m_2142_io_out_1)
  );
  Half_Adder m_2143 ( // @[MUL.scala 124:19]
    .io_in_0(m_2143_io_in_0),
    .io_in_1(m_2143_io_in_1),
    .io_out_0(m_2143_io_out_0),
    .io_out_1(m_2143_io_out_1)
  );
  Half_Adder m_2144 ( // @[MUL.scala 124:19]
    .io_in_0(m_2144_io_in_0),
    .io_in_1(m_2144_io_in_1),
    .io_out_0(m_2144_io_out_0),
    .io_out_1(m_2144_io_out_1)
  );
  Half_Adder m_2145 ( // @[MUL.scala 124:19]
    .io_in_0(m_2145_io_in_0),
    .io_in_1(m_2145_io_in_1),
    .io_out_0(m_2145_io_out_0),
    .io_out_1(m_2145_io_out_1)
  );
  Half_Adder m_2146 ( // @[MUL.scala 124:19]
    .io_in_0(m_2146_io_in_0),
    .io_in_1(m_2146_io_in_1),
    .io_out_0(m_2146_io_out_0),
    .io_out_1(m_2146_io_out_1)
  );
  Half_Adder m_2147 ( // @[MUL.scala 124:19]
    .io_in_0(m_2147_io_in_0),
    .io_in_1(m_2147_io_in_1),
    .io_out_0(m_2147_io_out_0),
    .io_out_1(m_2147_io_out_1)
  );
  Half_Adder m_2148 ( // @[MUL.scala 124:19]
    .io_in_0(m_2148_io_in_0),
    .io_in_1(m_2148_io_in_1),
    .io_out_0(m_2148_io_out_0),
    .io_out_1(m_2148_io_out_1)
  );
  Half_Adder m_2149 ( // @[MUL.scala 124:19]
    .io_in_0(m_2149_io_in_0),
    .io_in_1(m_2149_io_in_1),
    .io_out_0(m_2149_io_out_0),
    .io_out_1(m_2149_io_out_1)
  );
  Half_Adder m_2150 ( // @[MUL.scala 124:19]
    .io_in_0(m_2150_io_in_0),
    .io_in_1(m_2150_io_in_1),
    .io_out_0(m_2150_io_out_0),
    .io_out_1(m_2150_io_out_1)
  );
  Half_Adder m_2151 ( // @[MUL.scala 124:19]
    .io_in_0(m_2151_io_in_0),
    .io_in_1(m_2151_io_in_1),
    .io_out_0(m_2151_io_out_0),
    .io_out_1(m_2151_io_out_1)
  );
  Half_Adder m_2152 ( // @[MUL.scala 124:19]
    .io_in_0(m_2152_io_in_0),
    .io_in_1(m_2152_io_in_1),
    .io_out_0(m_2152_io_out_0),
    .io_out_1(m_2152_io_out_1)
  );
  Half_Adder m_2153 ( // @[MUL.scala 124:19]
    .io_in_0(m_2153_io_in_0),
    .io_in_1(m_2153_io_in_1),
    .io_out_0(m_2153_io_out_0),
    .io_out_1(m_2153_io_out_1)
  );
  Half_Adder m_2154 ( // @[MUL.scala 124:19]
    .io_in_0(m_2154_io_in_0),
    .io_in_1(m_2154_io_in_1),
    .io_out_0(m_2154_io_out_0),
    .io_out_1(m_2154_io_out_1)
  );
  Half_Adder m_2155 ( // @[MUL.scala 124:19]
    .io_in_0(m_2155_io_in_0),
    .io_in_1(m_2155_io_in_1),
    .io_out_0(m_2155_io_out_0),
    .io_out_1(m_2155_io_out_1)
  );
  Half_Adder m_2156 ( // @[MUL.scala 124:19]
    .io_in_0(m_2156_io_in_0),
    .io_in_1(m_2156_io_in_1),
    .io_out_0(m_2156_io_out_0),
    .io_out_1(m_2156_io_out_1)
  );
  Half_Adder m_2157 ( // @[MUL.scala 124:19]
    .io_in_0(m_2157_io_in_0),
    .io_in_1(m_2157_io_in_1),
    .io_out_0(m_2157_io_out_0),
    .io_out_1(m_2157_io_out_1)
  );
  Half_Adder m_2158 ( // @[MUL.scala 124:19]
    .io_in_0(m_2158_io_in_0),
    .io_in_1(m_2158_io_in_1),
    .io_out_0(m_2158_io_out_0),
    .io_out_1(m_2158_io_out_1)
  );
  Half_Adder m_2159 ( // @[MUL.scala 124:19]
    .io_in_0(m_2159_io_in_0),
    .io_in_1(m_2159_io_in_1),
    .io_out_0(m_2159_io_out_0),
    .io_out_1(m_2159_io_out_1)
  );
  Adder m_2160 ( // @[MUL.scala 102:19]
    .io_x1(m_2160_io_x1),
    .io_x2(m_2160_io_x2),
    .io_x3(m_2160_io_x3),
    .io_s(m_2160_io_s),
    .io_cout(m_2160_io_cout)
  );
  Adder m_2161 ( // @[MUL.scala 102:19]
    .io_x1(m_2161_io_x1),
    .io_x2(m_2161_io_x2),
    .io_x3(m_2161_io_x3),
    .io_s(m_2161_io_s),
    .io_cout(m_2161_io_cout)
  );
  Adder m_2162 ( // @[MUL.scala 102:19]
    .io_x1(m_2162_io_x1),
    .io_x2(m_2162_io_x2),
    .io_x3(m_2162_io_x3),
    .io_s(m_2162_io_s),
    .io_cout(m_2162_io_cout)
  );
  Adder m_2163 ( // @[MUL.scala 102:19]
    .io_x1(m_2163_io_x1),
    .io_x2(m_2163_io_x2),
    .io_x3(m_2163_io_x3),
    .io_s(m_2163_io_s),
    .io_cout(m_2163_io_cout)
  );
  Adder m_2164 ( // @[MUL.scala 102:19]
    .io_x1(m_2164_io_x1),
    .io_x2(m_2164_io_x2),
    .io_x3(m_2164_io_x3),
    .io_s(m_2164_io_s),
    .io_cout(m_2164_io_cout)
  );
  Adder m_2165 ( // @[MUL.scala 102:19]
    .io_x1(m_2165_io_x1),
    .io_x2(m_2165_io_x2),
    .io_x3(m_2165_io_x3),
    .io_s(m_2165_io_s),
    .io_cout(m_2165_io_cout)
  );
  Adder m_2166 ( // @[MUL.scala 102:19]
    .io_x1(m_2166_io_x1),
    .io_x2(m_2166_io_x2),
    .io_x3(m_2166_io_x3),
    .io_s(m_2166_io_s),
    .io_cout(m_2166_io_cout)
  );
  Adder m_2167 ( // @[MUL.scala 102:19]
    .io_x1(m_2167_io_x1),
    .io_x2(m_2167_io_x2),
    .io_x3(m_2167_io_x3),
    .io_s(m_2167_io_s),
    .io_cout(m_2167_io_cout)
  );
  Adder m_2168 ( // @[MUL.scala 102:19]
    .io_x1(m_2168_io_x1),
    .io_x2(m_2168_io_x2),
    .io_x3(m_2168_io_x3),
    .io_s(m_2168_io_s),
    .io_cout(m_2168_io_cout)
  );
  Adder m_2169 ( // @[MUL.scala 102:19]
    .io_x1(m_2169_io_x1),
    .io_x2(m_2169_io_x2),
    .io_x3(m_2169_io_x3),
    .io_s(m_2169_io_s),
    .io_cout(m_2169_io_cout)
  );
  Adder m_2170 ( // @[MUL.scala 102:19]
    .io_x1(m_2170_io_x1),
    .io_x2(m_2170_io_x2),
    .io_x3(m_2170_io_x3),
    .io_s(m_2170_io_s),
    .io_cout(m_2170_io_cout)
  );
  Adder m_2171 ( // @[MUL.scala 102:19]
    .io_x1(m_2171_io_x1),
    .io_x2(m_2171_io_x2),
    .io_x3(m_2171_io_x3),
    .io_s(m_2171_io_s),
    .io_cout(m_2171_io_cout)
  );
  Adder m_2172 ( // @[MUL.scala 102:19]
    .io_x1(m_2172_io_x1),
    .io_x2(m_2172_io_x2),
    .io_x3(m_2172_io_x3),
    .io_s(m_2172_io_s),
    .io_cout(m_2172_io_cout)
  );
  Adder m_2173 ( // @[MUL.scala 102:19]
    .io_x1(m_2173_io_x1),
    .io_x2(m_2173_io_x2),
    .io_x3(m_2173_io_x3),
    .io_s(m_2173_io_s),
    .io_cout(m_2173_io_cout)
  );
  Adder m_2174 ( // @[MUL.scala 102:19]
    .io_x1(m_2174_io_x1),
    .io_x2(m_2174_io_x2),
    .io_x3(m_2174_io_x3),
    .io_s(m_2174_io_s),
    .io_cout(m_2174_io_cout)
  );
  Adder m_2175 ( // @[MUL.scala 102:19]
    .io_x1(m_2175_io_x1),
    .io_x2(m_2175_io_x2),
    .io_x3(m_2175_io_x3),
    .io_s(m_2175_io_s),
    .io_cout(m_2175_io_cout)
  );
  Adder m_2176 ( // @[MUL.scala 102:19]
    .io_x1(m_2176_io_x1),
    .io_x2(m_2176_io_x2),
    .io_x3(m_2176_io_x3),
    .io_s(m_2176_io_s),
    .io_cout(m_2176_io_cout)
  );
  Adder m_2177 ( // @[MUL.scala 102:19]
    .io_x1(m_2177_io_x1),
    .io_x2(m_2177_io_x2),
    .io_x3(m_2177_io_x3),
    .io_s(m_2177_io_s),
    .io_cout(m_2177_io_cout)
  );
  Adder m_2178 ( // @[MUL.scala 102:19]
    .io_x1(m_2178_io_x1),
    .io_x2(m_2178_io_x2),
    .io_x3(m_2178_io_x3),
    .io_s(m_2178_io_s),
    .io_cout(m_2178_io_cout)
  );
  Adder m_2179 ( // @[MUL.scala 102:19]
    .io_x1(m_2179_io_x1),
    .io_x2(m_2179_io_x2),
    .io_x3(m_2179_io_x3),
    .io_s(m_2179_io_s),
    .io_cout(m_2179_io_cout)
  );
  Adder m_2180 ( // @[MUL.scala 102:19]
    .io_x1(m_2180_io_x1),
    .io_x2(m_2180_io_x2),
    .io_x3(m_2180_io_x3),
    .io_s(m_2180_io_s),
    .io_cout(m_2180_io_cout)
  );
  Adder m_2181 ( // @[MUL.scala 102:19]
    .io_x1(m_2181_io_x1),
    .io_x2(m_2181_io_x2),
    .io_x3(m_2181_io_x3),
    .io_s(m_2181_io_s),
    .io_cout(m_2181_io_cout)
  );
  Adder m_2182 ( // @[MUL.scala 102:19]
    .io_x1(m_2182_io_x1),
    .io_x2(m_2182_io_x2),
    .io_x3(m_2182_io_x3),
    .io_s(m_2182_io_s),
    .io_cout(m_2182_io_cout)
  );
  Adder m_2183 ( // @[MUL.scala 102:19]
    .io_x1(m_2183_io_x1),
    .io_x2(m_2183_io_x2),
    .io_x3(m_2183_io_x3),
    .io_s(m_2183_io_s),
    .io_cout(m_2183_io_cout)
  );
  Adder m_2184 ( // @[MUL.scala 102:19]
    .io_x1(m_2184_io_x1),
    .io_x2(m_2184_io_x2),
    .io_x3(m_2184_io_x3),
    .io_s(m_2184_io_s),
    .io_cout(m_2184_io_cout)
  );
  Adder m_2185 ( // @[MUL.scala 102:19]
    .io_x1(m_2185_io_x1),
    .io_x2(m_2185_io_x2),
    .io_x3(m_2185_io_x3),
    .io_s(m_2185_io_s),
    .io_cout(m_2185_io_cout)
  );
  Adder m_2186 ( // @[MUL.scala 102:19]
    .io_x1(m_2186_io_x1),
    .io_x2(m_2186_io_x2),
    .io_x3(m_2186_io_x3),
    .io_s(m_2186_io_s),
    .io_cout(m_2186_io_cout)
  );
  Adder m_2187 ( // @[MUL.scala 102:19]
    .io_x1(m_2187_io_x1),
    .io_x2(m_2187_io_x2),
    .io_x3(m_2187_io_x3),
    .io_s(m_2187_io_s),
    .io_cout(m_2187_io_cout)
  );
  Adder m_2188 ( // @[MUL.scala 102:19]
    .io_x1(m_2188_io_x1),
    .io_x2(m_2188_io_x2),
    .io_x3(m_2188_io_x3),
    .io_s(m_2188_io_s),
    .io_cout(m_2188_io_cout)
  );
  Adder m_2189 ( // @[MUL.scala 102:19]
    .io_x1(m_2189_io_x1),
    .io_x2(m_2189_io_x2),
    .io_x3(m_2189_io_x3),
    .io_s(m_2189_io_s),
    .io_cout(m_2189_io_cout)
  );
  Adder m_2190 ( // @[MUL.scala 102:19]
    .io_x1(m_2190_io_x1),
    .io_x2(m_2190_io_x2),
    .io_x3(m_2190_io_x3),
    .io_s(m_2190_io_s),
    .io_cout(m_2190_io_cout)
  );
  Adder m_2191 ( // @[MUL.scala 102:19]
    .io_x1(m_2191_io_x1),
    .io_x2(m_2191_io_x2),
    .io_x3(m_2191_io_x3),
    .io_s(m_2191_io_s),
    .io_cout(m_2191_io_cout)
  );
  Half_Adder m_2192 ( // @[MUL.scala 124:19]
    .io_in_0(m_2192_io_in_0),
    .io_in_1(m_2192_io_in_1),
    .io_out_0(m_2192_io_out_0),
    .io_out_1(m_2192_io_out_1)
  );
  Adder m_2193 ( // @[MUL.scala 102:19]
    .io_x1(m_2193_io_x1),
    .io_x2(m_2193_io_x2),
    .io_x3(m_2193_io_x3),
    .io_s(m_2193_io_s),
    .io_cout(m_2193_io_cout)
  );
  Half_Adder m_2194 ( // @[MUL.scala 124:19]
    .io_in_0(m_2194_io_in_0),
    .io_in_1(m_2194_io_in_1),
    .io_out_0(m_2194_io_out_0),
    .io_out_1(m_2194_io_out_1)
  );
  Adder m_2195 ( // @[MUL.scala 102:19]
    .io_x1(m_2195_io_x1),
    .io_x2(m_2195_io_x2),
    .io_x3(m_2195_io_x3),
    .io_s(m_2195_io_s),
    .io_cout(m_2195_io_cout)
  );
  Half_Adder m_2196 ( // @[MUL.scala 124:19]
    .io_in_0(m_2196_io_in_0),
    .io_in_1(m_2196_io_in_1),
    .io_out_0(m_2196_io_out_0),
    .io_out_1(m_2196_io_out_1)
  );
  Adder m_2197 ( // @[MUL.scala 102:19]
    .io_x1(m_2197_io_x1),
    .io_x2(m_2197_io_x2),
    .io_x3(m_2197_io_x3),
    .io_s(m_2197_io_s),
    .io_cout(m_2197_io_cout)
  );
  Half_Adder m_2198 ( // @[MUL.scala 124:19]
    .io_in_0(m_2198_io_in_0),
    .io_in_1(m_2198_io_in_1),
    .io_out_0(m_2198_io_out_0),
    .io_out_1(m_2198_io_out_1)
  );
  Adder m_2199 ( // @[MUL.scala 102:19]
    .io_x1(m_2199_io_x1),
    .io_x2(m_2199_io_x2),
    .io_x3(m_2199_io_x3),
    .io_s(m_2199_io_s),
    .io_cout(m_2199_io_cout)
  );
  Half_Adder m_2200 ( // @[MUL.scala 124:19]
    .io_in_0(m_2200_io_in_0),
    .io_in_1(m_2200_io_in_1),
    .io_out_0(m_2200_io_out_0),
    .io_out_1(m_2200_io_out_1)
  );
  Adder m_2201 ( // @[MUL.scala 102:19]
    .io_x1(m_2201_io_x1),
    .io_x2(m_2201_io_x2),
    .io_x3(m_2201_io_x3),
    .io_s(m_2201_io_s),
    .io_cout(m_2201_io_cout)
  );
  Half_Adder m_2202 ( // @[MUL.scala 124:19]
    .io_in_0(m_2202_io_in_0),
    .io_in_1(m_2202_io_in_1),
    .io_out_0(m_2202_io_out_0),
    .io_out_1(m_2202_io_out_1)
  );
  Adder m_2203 ( // @[MUL.scala 102:19]
    .io_x1(m_2203_io_x1),
    .io_x2(m_2203_io_x2),
    .io_x3(m_2203_io_x3),
    .io_s(m_2203_io_s),
    .io_cout(m_2203_io_cout)
  );
  Half_Adder m_2204 ( // @[MUL.scala 124:19]
    .io_in_0(m_2204_io_in_0),
    .io_in_1(m_2204_io_in_1),
    .io_out_0(m_2204_io_out_0),
    .io_out_1(m_2204_io_out_1)
  );
  Adder m_2205 ( // @[MUL.scala 102:19]
    .io_x1(m_2205_io_x1),
    .io_x2(m_2205_io_x2),
    .io_x3(m_2205_io_x3),
    .io_s(m_2205_io_s),
    .io_cout(m_2205_io_cout)
  );
  Half_Adder m_2206 ( // @[MUL.scala 124:19]
    .io_in_0(m_2206_io_in_0),
    .io_in_1(m_2206_io_in_1),
    .io_out_0(m_2206_io_out_0),
    .io_out_1(m_2206_io_out_1)
  );
  Adder m_2207 ( // @[MUL.scala 102:19]
    .io_x1(m_2207_io_x1),
    .io_x2(m_2207_io_x2),
    .io_x3(m_2207_io_x3),
    .io_s(m_2207_io_s),
    .io_cout(m_2207_io_cout)
  );
  Half_Adder m_2208 ( // @[MUL.scala 124:19]
    .io_in_0(m_2208_io_in_0),
    .io_in_1(m_2208_io_in_1),
    .io_out_0(m_2208_io_out_0),
    .io_out_1(m_2208_io_out_1)
  );
  Adder m_2209 ( // @[MUL.scala 102:19]
    .io_x1(m_2209_io_x1),
    .io_x2(m_2209_io_x2),
    .io_x3(m_2209_io_x3),
    .io_s(m_2209_io_s),
    .io_cout(m_2209_io_cout)
  );
  Half_Adder m_2210 ( // @[MUL.scala 124:19]
    .io_in_0(m_2210_io_in_0),
    .io_in_1(m_2210_io_in_1),
    .io_out_0(m_2210_io_out_0),
    .io_out_1(m_2210_io_out_1)
  );
  Adder m_2211 ( // @[MUL.scala 102:19]
    .io_x1(m_2211_io_x1),
    .io_x2(m_2211_io_x2),
    .io_x3(m_2211_io_x3),
    .io_s(m_2211_io_s),
    .io_cout(m_2211_io_cout)
  );
  Half_Adder m_2212 ( // @[MUL.scala 124:19]
    .io_in_0(m_2212_io_in_0),
    .io_in_1(m_2212_io_in_1),
    .io_out_0(m_2212_io_out_0),
    .io_out_1(m_2212_io_out_1)
  );
  Adder m_2213 ( // @[MUL.scala 102:19]
    .io_x1(m_2213_io_x1),
    .io_x2(m_2213_io_x2),
    .io_x3(m_2213_io_x3),
    .io_s(m_2213_io_s),
    .io_cout(m_2213_io_cout)
  );
  Half_Adder m_2214 ( // @[MUL.scala 124:19]
    .io_in_0(m_2214_io_in_0),
    .io_in_1(m_2214_io_in_1),
    .io_out_0(m_2214_io_out_0),
    .io_out_1(m_2214_io_out_1)
  );
  Adder m_2215 ( // @[MUL.scala 102:19]
    .io_x1(m_2215_io_x1),
    .io_x2(m_2215_io_x2),
    .io_x3(m_2215_io_x3),
    .io_s(m_2215_io_s),
    .io_cout(m_2215_io_cout)
  );
  Half_Adder m_2216 ( // @[MUL.scala 124:19]
    .io_in_0(m_2216_io_in_0),
    .io_in_1(m_2216_io_in_1),
    .io_out_0(m_2216_io_out_0),
    .io_out_1(m_2216_io_out_1)
  );
  Adder m_2217 ( // @[MUL.scala 102:19]
    .io_x1(m_2217_io_x1),
    .io_x2(m_2217_io_x2),
    .io_x3(m_2217_io_x3),
    .io_s(m_2217_io_s),
    .io_cout(m_2217_io_cout)
  );
  Half_Adder m_2218 ( // @[MUL.scala 124:19]
    .io_in_0(m_2218_io_in_0),
    .io_in_1(m_2218_io_in_1),
    .io_out_0(m_2218_io_out_0),
    .io_out_1(m_2218_io_out_1)
  );
  Adder m_2219 ( // @[MUL.scala 102:19]
    .io_x1(m_2219_io_x1),
    .io_x2(m_2219_io_x2),
    .io_x3(m_2219_io_x3),
    .io_s(m_2219_io_s),
    .io_cout(m_2219_io_cout)
  );
  Half_Adder m_2220 ( // @[MUL.scala 124:19]
    .io_in_0(m_2220_io_in_0),
    .io_in_1(m_2220_io_in_1),
    .io_out_0(m_2220_io_out_0),
    .io_out_1(m_2220_io_out_1)
  );
  Adder m_2221 ( // @[MUL.scala 102:19]
    .io_x1(m_2221_io_x1),
    .io_x2(m_2221_io_x2),
    .io_x3(m_2221_io_x3),
    .io_s(m_2221_io_s),
    .io_cout(m_2221_io_cout)
  );
  Half_Adder m_2222 ( // @[MUL.scala 124:19]
    .io_in_0(m_2222_io_in_0),
    .io_in_1(m_2222_io_in_1),
    .io_out_0(m_2222_io_out_0),
    .io_out_1(m_2222_io_out_1)
  );
  Adder m_2223 ( // @[MUL.scala 102:19]
    .io_x1(m_2223_io_x1),
    .io_x2(m_2223_io_x2),
    .io_x3(m_2223_io_x3),
    .io_s(m_2223_io_s),
    .io_cout(m_2223_io_cout)
  );
  Half_Adder m_2224 ( // @[MUL.scala 124:19]
    .io_in_0(m_2224_io_in_0),
    .io_in_1(m_2224_io_in_1),
    .io_out_0(m_2224_io_out_0),
    .io_out_1(m_2224_io_out_1)
  );
  Adder m_2225 ( // @[MUL.scala 102:19]
    .io_x1(m_2225_io_x1),
    .io_x2(m_2225_io_x2),
    .io_x3(m_2225_io_x3),
    .io_s(m_2225_io_s),
    .io_cout(m_2225_io_cout)
  );
  Half_Adder m_2226 ( // @[MUL.scala 124:19]
    .io_in_0(m_2226_io_in_0),
    .io_in_1(m_2226_io_in_1),
    .io_out_0(m_2226_io_out_0),
    .io_out_1(m_2226_io_out_1)
  );
  Adder m_2227 ( // @[MUL.scala 102:19]
    .io_x1(m_2227_io_x1),
    .io_x2(m_2227_io_x2),
    .io_x3(m_2227_io_x3),
    .io_s(m_2227_io_s),
    .io_cout(m_2227_io_cout)
  );
  Half_Adder m_2228 ( // @[MUL.scala 124:19]
    .io_in_0(m_2228_io_in_0),
    .io_in_1(m_2228_io_in_1),
    .io_out_0(m_2228_io_out_0),
    .io_out_1(m_2228_io_out_1)
  );
  Adder m_2229 ( // @[MUL.scala 102:19]
    .io_x1(m_2229_io_x1),
    .io_x2(m_2229_io_x2),
    .io_x3(m_2229_io_x3),
    .io_s(m_2229_io_s),
    .io_cout(m_2229_io_cout)
  );
  Half_Adder m_2230 ( // @[MUL.scala 124:19]
    .io_in_0(m_2230_io_in_0),
    .io_in_1(m_2230_io_in_1),
    .io_out_0(m_2230_io_out_0),
    .io_out_1(m_2230_io_out_1)
  );
  Adder m_2231 ( // @[MUL.scala 102:19]
    .io_x1(m_2231_io_x1),
    .io_x2(m_2231_io_x2),
    .io_x3(m_2231_io_x3),
    .io_s(m_2231_io_s),
    .io_cout(m_2231_io_cout)
  );
  Half_Adder m_2232 ( // @[MUL.scala 124:19]
    .io_in_0(m_2232_io_in_0),
    .io_in_1(m_2232_io_in_1),
    .io_out_0(m_2232_io_out_0),
    .io_out_1(m_2232_io_out_1)
  );
  Adder m_2233 ( // @[MUL.scala 102:19]
    .io_x1(m_2233_io_x1),
    .io_x2(m_2233_io_x2),
    .io_x3(m_2233_io_x3),
    .io_s(m_2233_io_s),
    .io_cout(m_2233_io_cout)
  );
  Adder m_2234 ( // @[MUL.scala 102:19]
    .io_x1(m_2234_io_x1),
    .io_x2(m_2234_io_x2),
    .io_x3(m_2234_io_x3),
    .io_s(m_2234_io_s),
    .io_cout(m_2234_io_cout)
  );
  Adder m_2235 ( // @[MUL.scala 102:19]
    .io_x1(m_2235_io_x1),
    .io_x2(m_2235_io_x2),
    .io_x3(m_2235_io_x3),
    .io_s(m_2235_io_s),
    .io_cout(m_2235_io_cout)
  );
  Adder m_2236 ( // @[MUL.scala 102:19]
    .io_x1(m_2236_io_x1),
    .io_x2(m_2236_io_x2),
    .io_x3(m_2236_io_x3),
    .io_s(m_2236_io_s),
    .io_cout(m_2236_io_cout)
  );
  Adder m_2237 ( // @[MUL.scala 102:19]
    .io_x1(m_2237_io_x1),
    .io_x2(m_2237_io_x2),
    .io_x3(m_2237_io_x3),
    .io_s(m_2237_io_s),
    .io_cout(m_2237_io_cout)
  );
  Adder m_2238 ( // @[MUL.scala 102:19]
    .io_x1(m_2238_io_x1),
    .io_x2(m_2238_io_x2),
    .io_x3(m_2238_io_x3),
    .io_s(m_2238_io_s),
    .io_cout(m_2238_io_cout)
  );
  Adder m_2239 ( // @[MUL.scala 102:19]
    .io_x1(m_2239_io_x1),
    .io_x2(m_2239_io_x2),
    .io_x3(m_2239_io_x3),
    .io_s(m_2239_io_s),
    .io_cout(m_2239_io_cout)
  );
  Adder m_2240 ( // @[MUL.scala 102:19]
    .io_x1(m_2240_io_x1),
    .io_x2(m_2240_io_x2),
    .io_x3(m_2240_io_x3),
    .io_s(m_2240_io_s),
    .io_cout(m_2240_io_cout)
  );
  Adder m_2241 ( // @[MUL.scala 102:19]
    .io_x1(m_2241_io_x1),
    .io_x2(m_2241_io_x2),
    .io_x3(m_2241_io_x3),
    .io_s(m_2241_io_s),
    .io_cout(m_2241_io_cout)
  );
  Adder m_2242 ( // @[MUL.scala 102:19]
    .io_x1(m_2242_io_x1),
    .io_x2(m_2242_io_x2),
    .io_x3(m_2242_io_x3),
    .io_s(m_2242_io_s),
    .io_cout(m_2242_io_cout)
  );
  Adder m_2243 ( // @[MUL.scala 102:19]
    .io_x1(m_2243_io_x1),
    .io_x2(m_2243_io_x2),
    .io_x3(m_2243_io_x3),
    .io_s(m_2243_io_s),
    .io_cout(m_2243_io_cout)
  );
  Adder m_2244 ( // @[MUL.scala 102:19]
    .io_x1(m_2244_io_x1),
    .io_x2(m_2244_io_x2),
    .io_x3(m_2244_io_x3),
    .io_s(m_2244_io_s),
    .io_cout(m_2244_io_cout)
  );
  Adder m_2245 ( // @[MUL.scala 102:19]
    .io_x1(m_2245_io_x1),
    .io_x2(m_2245_io_x2),
    .io_x3(m_2245_io_x3),
    .io_s(m_2245_io_s),
    .io_cout(m_2245_io_cout)
  );
  Adder m_2246 ( // @[MUL.scala 102:19]
    .io_x1(m_2246_io_x1),
    .io_x2(m_2246_io_x2),
    .io_x3(m_2246_io_x3),
    .io_s(m_2246_io_s),
    .io_cout(m_2246_io_cout)
  );
  Adder m_2247 ( // @[MUL.scala 102:19]
    .io_x1(m_2247_io_x1),
    .io_x2(m_2247_io_x2),
    .io_x3(m_2247_io_x3),
    .io_s(m_2247_io_s),
    .io_cout(m_2247_io_cout)
  );
  Adder m_2248 ( // @[MUL.scala 102:19]
    .io_x1(m_2248_io_x1),
    .io_x2(m_2248_io_x2),
    .io_x3(m_2248_io_x3),
    .io_s(m_2248_io_s),
    .io_cout(m_2248_io_cout)
  );
  Adder m_2249 ( // @[MUL.scala 102:19]
    .io_x1(m_2249_io_x1),
    .io_x2(m_2249_io_x2),
    .io_x3(m_2249_io_x3),
    .io_s(m_2249_io_s),
    .io_cout(m_2249_io_cout)
  );
  Adder m_2250 ( // @[MUL.scala 102:19]
    .io_x1(m_2250_io_x1),
    .io_x2(m_2250_io_x2),
    .io_x3(m_2250_io_x3),
    .io_s(m_2250_io_s),
    .io_cout(m_2250_io_cout)
  );
  Adder m_2251 ( // @[MUL.scala 102:19]
    .io_x1(m_2251_io_x1),
    .io_x2(m_2251_io_x2),
    .io_x3(m_2251_io_x3),
    .io_s(m_2251_io_s),
    .io_cout(m_2251_io_cout)
  );
  Adder m_2252 ( // @[MUL.scala 102:19]
    .io_x1(m_2252_io_x1),
    .io_x2(m_2252_io_x2),
    .io_x3(m_2252_io_x3),
    .io_s(m_2252_io_s),
    .io_cout(m_2252_io_cout)
  );
  Adder m_2253 ( // @[MUL.scala 102:19]
    .io_x1(m_2253_io_x1),
    .io_x2(m_2253_io_x2),
    .io_x3(m_2253_io_x3),
    .io_s(m_2253_io_s),
    .io_cout(m_2253_io_cout)
  );
  Adder m_2254 ( // @[MUL.scala 102:19]
    .io_x1(m_2254_io_x1),
    .io_x2(m_2254_io_x2),
    .io_x3(m_2254_io_x3),
    .io_s(m_2254_io_s),
    .io_cout(m_2254_io_cout)
  );
  Adder m_2255 ( // @[MUL.scala 102:19]
    .io_x1(m_2255_io_x1),
    .io_x2(m_2255_io_x2),
    .io_x3(m_2255_io_x3),
    .io_s(m_2255_io_s),
    .io_cout(m_2255_io_cout)
  );
  Adder m_2256 ( // @[MUL.scala 102:19]
    .io_x1(m_2256_io_x1),
    .io_x2(m_2256_io_x2),
    .io_x3(m_2256_io_x3),
    .io_s(m_2256_io_s),
    .io_cout(m_2256_io_cout)
  );
  Adder m_2257 ( // @[MUL.scala 102:19]
    .io_x1(m_2257_io_x1),
    .io_x2(m_2257_io_x2),
    .io_x3(m_2257_io_x3),
    .io_s(m_2257_io_s),
    .io_cout(m_2257_io_cout)
  );
  Adder m_2258 ( // @[MUL.scala 102:19]
    .io_x1(m_2258_io_x1),
    .io_x2(m_2258_io_x2),
    .io_x3(m_2258_io_x3),
    .io_s(m_2258_io_s),
    .io_cout(m_2258_io_cout)
  );
  Adder m_2259 ( // @[MUL.scala 102:19]
    .io_x1(m_2259_io_x1),
    .io_x2(m_2259_io_x2),
    .io_x3(m_2259_io_x3),
    .io_s(m_2259_io_s),
    .io_cout(m_2259_io_cout)
  );
  Adder m_2260 ( // @[MUL.scala 102:19]
    .io_x1(m_2260_io_x1),
    .io_x2(m_2260_io_x2),
    .io_x3(m_2260_io_x3),
    .io_s(m_2260_io_s),
    .io_cout(m_2260_io_cout)
  );
  Adder m_2261 ( // @[MUL.scala 102:19]
    .io_x1(m_2261_io_x1),
    .io_x2(m_2261_io_x2),
    .io_x3(m_2261_io_x3),
    .io_s(m_2261_io_s),
    .io_cout(m_2261_io_cout)
  );
  Adder m_2262 ( // @[MUL.scala 102:19]
    .io_x1(m_2262_io_x1),
    .io_x2(m_2262_io_x2),
    .io_x3(m_2262_io_x3),
    .io_s(m_2262_io_s),
    .io_cout(m_2262_io_cout)
  );
  Half_Adder m_2263 ( // @[MUL.scala 124:19]
    .io_in_0(m_2263_io_in_0),
    .io_in_1(m_2263_io_in_1),
    .io_out_0(m_2263_io_out_0),
    .io_out_1(m_2263_io_out_1)
  );
  Half_Adder m_2264 ( // @[MUL.scala 124:19]
    .io_in_0(m_2264_io_in_0),
    .io_in_1(m_2264_io_in_1),
    .io_out_0(m_2264_io_out_0),
    .io_out_1(m_2264_io_out_1)
  );
  Half_Adder m_2265 ( // @[MUL.scala 124:19]
    .io_in_0(m_2265_io_in_0),
    .io_in_1(m_2265_io_in_1),
    .io_out_0(m_2265_io_out_0),
    .io_out_1(m_2265_io_out_1)
  );
  Half_Adder m_2266 ( // @[MUL.scala 124:19]
    .io_in_0(m_2266_io_in_0),
    .io_in_1(m_2266_io_in_1),
    .io_out_0(m_2266_io_out_0),
    .io_out_1(m_2266_io_out_1)
  );
  Half_Adder m_2267 ( // @[MUL.scala 124:19]
    .io_in_0(m_2267_io_in_0),
    .io_in_1(m_2267_io_in_1),
    .io_out_0(m_2267_io_out_0),
    .io_out_1(m_2267_io_out_1)
  );
  Half_Adder m_2268 ( // @[MUL.scala 124:19]
    .io_in_0(m_2268_io_in_0),
    .io_in_1(m_2268_io_in_1),
    .io_out_0(m_2268_io_out_0),
    .io_out_1(m_2268_io_out_1)
  );
  Half_Adder m_2269 ( // @[MUL.scala 124:19]
    .io_in_0(m_2269_io_in_0),
    .io_in_1(m_2269_io_in_1),
    .io_out_0(m_2269_io_out_0),
    .io_out_1(m_2269_io_out_1)
  );
  Half_Adder m_2270 ( // @[MUL.scala 124:19]
    .io_in_0(m_2270_io_in_0),
    .io_in_1(m_2270_io_in_1),
    .io_out_0(m_2270_io_out_0),
    .io_out_1(m_2270_io_out_1)
  );
  Half_Adder m_2271 ( // @[MUL.scala 124:19]
    .io_in_0(m_2271_io_in_0),
    .io_in_1(m_2271_io_in_1),
    .io_out_0(m_2271_io_out_0),
    .io_out_1(m_2271_io_out_1)
  );
  Half_Adder m_2272 ( // @[MUL.scala 124:19]
    .io_in_0(m_2272_io_in_0),
    .io_in_1(m_2272_io_in_1),
    .io_out_0(m_2272_io_out_0),
    .io_out_1(m_2272_io_out_1)
  );
  Half_Adder m_2273 ( // @[MUL.scala 124:19]
    .io_in_0(m_2273_io_in_0),
    .io_in_1(m_2273_io_in_1),
    .io_out_0(m_2273_io_out_0),
    .io_out_1(m_2273_io_out_1)
  );
  Half_Adder m_2274 ( // @[MUL.scala 124:19]
    .io_in_0(m_2274_io_in_0),
    .io_in_1(m_2274_io_in_1),
    .io_out_0(m_2274_io_out_0),
    .io_out_1(m_2274_io_out_1)
  );
  Half_Adder m_2275 ( // @[MUL.scala 124:19]
    .io_in_0(m_2275_io_in_0),
    .io_in_1(m_2275_io_in_1),
    .io_out_0(m_2275_io_out_0),
    .io_out_1(m_2275_io_out_1)
  );
  Half_Adder m_2276 ( // @[MUL.scala 124:19]
    .io_in_0(m_2276_io_in_0),
    .io_in_1(m_2276_io_in_1),
    .io_out_0(m_2276_io_out_0),
    .io_out_1(m_2276_io_out_1)
  );
  Half_Adder m_2277 ( // @[MUL.scala 124:19]
    .io_in_0(m_2277_io_in_0),
    .io_in_1(m_2277_io_in_1),
    .io_out_0(m_2277_io_out_0),
    .io_out_1(m_2277_io_out_1)
  );
  Half_Adder m_2278 ( // @[MUL.scala 124:19]
    .io_in_0(m_2278_io_in_0),
    .io_in_1(m_2278_io_in_1),
    .io_out_0(m_2278_io_out_0),
    .io_out_1(m_2278_io_out_1)
  );
  Half_Adder m_2279 ( // @[MUL.scala 124:19]
    .io_in_0(m_2279_io_in_0),
    .io_in_1(m_2279_io_in_1),
    .io_out_0(m_2279_io_out_0),
    .io_out_1(m_2279_io_out_1)
  );
  Half_Adder m_2280 ( // @[MUL.scala 124:19]
    .io_in_0(m_2280_io_in_0),
    .io_in_1(m_2280_io_in_1),
    .io_out_0(m_2280_io_out_0),
    .io_out_1(m_2280_io_out_1)
  );
  Half_Adder m_2281 ( // @[MUL.scala 124:19]
    .io_in_0(m_2281_io_in_0),
    .io_in_1(m_2281_io_in_1),
    .io_out_0(m_2281_io_out_0),
    .io_out_1(m_2281_io_out_1)
  );
  Half_Adder m_2282 ( // @[MUL.scala 124:19]
    .io_in_0(m_2282_io_in_0),
    .io_in_1(m_2282_io_in_1),
    .io_out_0(m_2282_io_out_0),
    .io_out_1(m_2282_io_out_1)
  );
  Half_Adder m_2283 ( // @[MUL.scala 124:19]
    .io_in_0(m_2283_io_in_0),
    .io_in_1(m_2283_io_in_1),
    .io_out_0(m_2283_io_out_0),
    .io_out_1(m_2283_io_out_1)
  );
  Half_Adder m_2284 ( // @[MUL.scala 124:19]
    .io_in_0(m_2284_io_in_0),
    .io_in_1(m_2284_io_in_1),
    .io_out_0(m_2284_io_out_0),
    .io_out_1(m_2284_io_out_1)
  );
  Half_Adder m_2285 ( // @[MUL.scala 124:19]
    .io_in_0(m_2285_io_in_0),
    .io_in_1(m_2285_io_in_1),
    .io_out_0(m_2285_io_out_0),
    .io_out_1(m_2285_io_out_1)
  );
  Half_Adder m_2286 ( // @[MUL.scala 124:19]
    .io_in_0(m_2286_io_in_0),
    .io_in_1(m_2286_io_in_1),
    .io_out_0(m_2286_io_out_0),
    .io_out_1(m_2286_io_out_1)
  );
  Half_Adder m_2287 ( // @[MUL.scala 124:19]
    .io_in_0(m_2287_io_in_0),
    .io_in_1(m_2287_io_in_1),
    .io_out_0(m_2287_io_out_0),
    .io_out_1(m_2287_io_out_1)
  );
  Half_Adder m_2288 ( // @[MUL.scala 124:19]
    .io_in_0(m_2288_io_in_0),
    .io_in_1(m_2288_io_in_1),
    .io_out_0(m_2288_io_out_0),
    .io_out_1(m_2288_io_out_1)
  );
  Half_Adder m_2289 ( // @[MUL.scala 124:19]
    .io_in_0(m_2289_io_in_0),
    .io_in_1(m_2289_io_in_1),
    .io_out_0(m_2289_io_out_0),
    .io_out_1(m_2289_io_out_1)
  );
  Half_Adder m_2290 ( // @[MUL.scala 124:19]
    .io_in_0(m_2290_io_in_0),
    .io_in_1(m_2290_io_in_1),
    .io_out_0(m_2290_io_out_0),
    .io_out_1(m_2290_io_out_1)
  );
  Half_Adder m_2291 ( // @[MUL.scala 124:19]
    .io_in_0(m_2291_io_in_0),
    .io_in_1(m_2291_io_in_1),
    .io_out_0(m_2291_io_out_0),
    .io_out_1(m_2291_io_out_1)
  );
  Half_Adder m_2292 ( // @[MUL.scala 124:19]
    .io_in_0(m_2292_io_in_0),
    .io_in_1(m_2292_io_in_1),
    .io_out_0(m_2292_io_out_0),
    .io_out_1(m_2292_io_out_1)
  );
  Half_Adder m_2293 ( // @[MUL.scala 124:19]
    .io_in_0(m_2293_io_in_0),
    .io_in_1(m_2293_io_in_1),
    .io_out_0(m_2293_io_out_0),
    .io_out_1(m_2293_io_out_1)
  );
  Half_Adder m_2294 ( // @[MUL.scala 124:19]
    .io_in_0(m_2294_io_in_0),
    .io_in_1(m_2294_io_in_1),
    .io_out_0(m_2294_io_out_0),
    .io_out_1(m_2294_io_out_1)
  );
  Half_Adder m_2295 ( // @[MUL.scala 124:19]
    .io_in_0(m_2295_io_in_0),
    .io_in_1(m_2295_io_in_1),
    .io_out_0(m_2295_io_out_0),
    .io_out_1(m_2295_io_out_1)
  );
  Half_Adder m_2296 ( // @[MUL.scala 124:19]
    .io_in_0(m_2296_io_in_0),
    .io_in_1(m_2296_io_in_1),
    .io_out_0(m_2296_io_out_0),
    .io_out_1(m_2296_io_out_1)
  );
  Half_Adder m_2297 ( // @[MUL.scala 124:19]
    .io_in_0(m_2297_io_in_0),
    .io_in_1(m_2297_io_in_1),
    .io_out_0(m_2297_io_out_0),
    .io_out_1(m_2297_io_out_1)
  );
  Half_Adder m_2298 ( // @[MUL.scala 124:19]
    .io_in_0(m_2298_io_in_0),
    .io_in_1(m_2298_io_in_1),
    .io_out_0(m_2298_io_out_0),
    .io_out_1(m_2298_io_out_1)
  );
  Half_Adder m_2299 ( // @[MUL.scala 124:19]
    .io_in_0(m_2299_io_in_0),
    .io_in_1(m_2299_io_in_1),
    .io_out_0(m_2299_io_out_0),
    .io_out_1(m_2299_io_out_1)
  );
  Half_Adder m_2300 ( // @[MUL.scala 124:19]
    .io_in_0(m_2300_io_in_0),
    .io_in_1(m_2300_io_in_1),
    .io_out_0(m_2300_io_out_0),
    .io_out_1(m_2300_io_out_1)
  );
  Half_Adder m_2301 ( // @[MUL.scala 124:19]
    .io_in_0(m_2301_io_in_0),
    .io_in_1(m_2301_io_in_1),
    .io_out_0(m_2301_io_out_0),
    .io_out_1(m_2301_io_out_1)
  );
  Half_Adder m_2302 ( // @[MUL.scala 124:19]
    .io_in_0(m_2302_io_in_0),
    .io_in_1(m_2302_io_in_1),
    .io_out_0(m_2302_io_out_0),
    .io_out_1(m_2302_io_out_1)
  );
  Half_Adder m_2303 ( // @[MUL.scala 124:19]
    .io_in_0(m_2303_io_in_0),
    .io_in_1(m_2303_io_in_1),
    .io_out_0(m_2303_io_out_0),
    .io_out_1(m_2303_io_out_1)
  );
  Half_Adder m_2304 ( // @[MUL.scala 124:19]
    .io_in_0(m_2304_io_in_0),
    .io_in_1(m_2304_io_in_1),
    .io_out_0(m_2304_io_out_0),
    .io_out_1(m_2304_io_out_1)
  );
  Half_Adder m_2305 ( // @[MUL.scala 124:19]
    .io_in_0(m_2305_io_in_0),
    .io_in_1(m_2305_io_in_1),
    .io_out_0(m_2305_io_out_0),
    .io_out_1(m_2305_io_out_1)
  );
  Half_Adder m_2306 ( // @[MUL.scala 124:19]
    .io_in_0(m_2306_io_in_0),
    .io_in_1(m_2306_io_in_1),
    .io_out_0(m_2306_io_out_0),
    .io_out_1(m_2306_io_out_1)
  );
  Half_Adder m_2307 ( // @[MUL.scala 124:19]
    .io_in_0(m_2307_io_in_0),
    .io_in_1(m_2307_io_in_1),
    .io_out_0(m_2307_io_out_0),
    .io_out_1(m_2307_io_out_1)
  );
  Half_Adder m_2308 ( // @[MUL.scala 124:19]
    .io_in_0(m_2308_io_in_0),
    .io_in_1(m_2308_io_in_1),
    .io_out_0(m_2308_io_out_0),
    .io_out_1(m_2308_io_out_1)
  );
  Half_Adder m_2309 ( // @[MUL.scala 124:19]
    .io_in_0(m_2309_io_in_0),
    .io_in_1(m_2309_io_in_1),
    .io_out_0(m_2309_io_out_0),
    .io_out_1(m_2309_io_out_1)
  );
  Half_Adder m_2310 ( // @[MUL.scala 124:19]
    .io_in_0(m_2310_io_in_0),
    .io_in_1(m_2310_io_in_1),
    .io_out_0(m_2310_io_out_0),
    .io_out_1(m_2310_io_out_1)
  );
  Half_Adder m_2311 ( // @[MUL.scala 124:19]
    .io_in_0(m_2311_io_in_0),
    .io_in_1(m_2311_io_in_1),
    .io_out_0(m_2311_io_out_0),
    .io_out_1(m_2311_io_out_1)
  );
  Half_Adder m_2312 ( // @[MUL.scala 124:19]
    .io_in_0(m_2312_io_in_0),
    .io_in_1(m_2312_io_in_1),
    .io_out_0(m_2312_io_out_0),
    .io_out_1(m_2312_io_out_1)
  );
  Half_Adder m_2313 ( // @[MUL.scala 124:19]
    .io_in_0(m_2313_io_in_0),
    .io_in_1(m_2313_io_in_1),
    .io_out_0(m_2313_io_out_0),
    .io_out_1(m_2313_io_out_1)
  );
  Half_Adder m_2314 ( // @[MUL.scala 124:19]
    .io_in_0(m_2314_io_in_0),
    .io_in_1(m_2314_io_in_1),
    .io_out_0(m_2314_io_out_0),
    .io_out_1(m_2314_io_out_1)
  );
  Half_Adder m_2315 ( // @[MUL.scala 124:19]
    .io_in_0(m_2315_io_in_0),
    .io_in_1(m_2315_io_in_1),
    .io_out_0(m_2315_io_out_0),
    .io_out_1(m_2315_io_out_1)
  );
  Half_Adder m_2316 ( // @[MUL.scala 124:19]
    .io_in_0(m_2316_io_in_0),
    .io_in_1(m_2316_io_in_1),
    .io_out_0(m_2316_io_out_0),
    .io_out_1(m_2316_io_out_1)
  );
  Half_Adder m_2317 ( // @[MUL.scala 124:19]
    .io_in_0(m_2317_io_in_0),
    .io_in_1(m_2317_io_in_1),
    .io_out_0(m_2317_io_out_0),
    .io_out_1(m_2317_io_out_1)
  );
  Half_Adder m_2318 ( // @[MUL.scala 124:19]
    .io_in_0(m_2318_io_in_0),
    .io_in_1(m_2318_io_in_1),
    .io_out_0(m_2318_io_out_0),
    .io_out_1(m_2318_io_out_1)
  );
  Adder m_2319 ( // @[MUL.scala 102:19]
    .io_x1(m_2319_io_x1),
    .io_x2(m_2319_io_x2),
    .io_x3(m_2319_io_x3),
    .io_s(m_2319_io_s),
    .io_cout(m_2319_io_cout)
  );
  Adder m_2320 ( // @[MUL.scala 102:19]
    .io_x1(m_2320_io_x1),
    .io_x2(m_2320_io_x2),
    .io_x3(m_2320_io_x3),
    .io_s(m_2320_io_s),
    .io_cout(m_2320_io_cout)
  );
  Adder m_2321 ( // @[MUL.scala 102:19]
    .io_x1(m_2321_io_x1),
    .io_x2(m_2321_io_x2),
    .io_x3(m_2321_io_x3),
    .io_s(m_2321_io_s),
    .io_cout(m_2321_io_cout)
  );
  Adder m_2322 ( // @[MUL.scala 102:19]
    .io_x1(m_2322_io_x1),
    .io_x2(m_2322_io_x2),
    .io_x3(m_2322_io_x3),
    .io_s(m_2322_io_s),
    .io_cout(m_2322_io_cout)
  );
  Adder m_2323 ( // @[MUL.scala 102:19]
    .io_x1(m_2323_io_x1),
    .io_x2(m_2323_io_x2),
    .io_x3(m_2323_io_x3),
    .io_s(m_2323_io_s),
    .io_cout(m_2323_io_cout)
  );
  Adder m_2324 ( // @[MUL.scala 102:19]
    .io_x1(m_2324_io_x1),
    .io_x2(m_2324_io_x2),
    .io_x3(m_2324_io_x3),
    .io_s(m_2324_io_s),
    .io_cout(m_2324_io_cout)
  );
  Adder m_2325 ( // @[MUL.scala 102:19]
    .io_x1(m_2325_io_x1),
    .io_x2(m_2325_io_x2),
    .io_x3(m_2325_io_x3),
    .io_s(m_2325_io_s),
    .io_cout(m_2325_io_cout)
  );
  Adder m_2326 ( // @[MUL.scala 102:19]
    .io_x1(m_2326_io_x1),
    .io_x2(m_2326_io_x2),
    .io_x3(m_2326_io_x3),
    .io_s(m_2326_io_s),
    .io_cout(m_2326_io_cout)
  );
  Adder m_2327 ( // @[MUL.scala 102:19]
    .io_x1(m_2327_io_x1),
    .io_x2(m_2327_io_x2),
    .io_x3(m_2327_io_x3),
    .io_s(m_2327_io_s),
    .io_cout(m_2327_io_cout)
  );
  Adder m_2328 ( // @[MUL.scala 102:19]
    .io_x1(m_2328_io_x1),
    .io_x2(m_2328_io_x2),
    .io_x3(m_2328_io_x3),
    .io_s(m_2328_io_s),
    .io_cout(m_2328_io_cout)
  );
  Adder m_2329 ( // @[MUL.scala 102:19]
    .io_x1(m_2329_io_x1),
    .io_x2(m_2329_io_x2),
    .io_x3(m_2329_io_x3),
    .io_s(m_2329_io_s),
    .io_cout(m_2329_io_cout)
  );
  Adder m_2330 ( // @[MUL.scala 102:19]
    .io_x1(m_2330_io_x1),
    .io_x2(m_2330_io_x2),
    .io_x3(m_2330_io_x3),
    .io_s(m_2330_io_s),
    .io_cout(m_2330_io_cout)
  );
  Adder m_2331 ( // @[MUL.scala 102:19]
    .io_x1(m_2331_io_x1),
    .io_x2(m_2331_io_x2),
    .io_x3(m_2331_io_x3),
    .io_s(m_2331_io_s),
    .io_cout(m_2331_io_cout)
  );
  Adder m_2332 ( // @[MUL.scala 102:19]
    .io_x1(m_2332_io_x1),
    .io_x2(m_2332_io_x2),
    .io_x3(m_2332_io_x3),
    .io_s(m_2332_io_s),
    .io_cout(m_2332_io_cout)
  );
  Adder m_2333 ( // @[MUL.scala 102:19]
    .io_x1(m_2333_io_x1),
    .io_x2(m_2333_io_x2),
    .io_x3(m_2333_io_x3),
    .io_s(m_2333_io_s),
    .io_cout(m_2333_io_cout)
  );
  Adder m_2334 ( // @[MUL.scala 102:19]
    .io_x1(m_2334_io_x1),
    .io_x2(m_2334_io_x2),
    .io_x3(m_2334_io_x3),
    .io_s(m_2334_io_s),
    .io_cout(m_2334_io_cout)
  );
  Adder m_2335 ( // @[MUL.scala 102:19]
    .io_x1(m_2335_io_x1),
    .io_x2(m_2335_io_x2),
    .io_x3(m_2335_io_x3),
    .io_s(m_2335_io_s),
    .io_cout(m_2335_io_cout)
  );
  Adder m_2336 ( // @[MUL.scala 102:19]
    .io_x1(m_2336_io_x1),
    .io_x2(m_2336_io_x2),
    .io_x3(m_2336_io_x3),
    .io_s(m_2336_io_s),
    .io_cout(m_2336_io_cout)
  );
  Adder m_2337 ( // @[MUL.scala 102:19]
    .io_x1(m_2337_io_x1),
    .io_x2(m_2337_io_x2),
    .io_x3(m_2337_io_x3),
    .io_s(m_2337_io_s),
    .io_cout(m_2337_io_cout)
  );
  Adder m_2338 ( // @[MUL.scala 102:19]
    .io_x1(m_2338_io_x1),
    .io_x2(m_2338_io_x2),
    .io_x3(m_2338_io_x3),
    .io_s(m_2338_io_s),
    .io_cout(m_2338_io_cout)
  );
  Adder m_2339 ( // @[MUL.scala 102:19]
    .io_x1(m_2339_io_x1),
    .io_x2(m_2339_io_x2),
    .io_x3(m_2339_io_x3),
    .io_s(m_2339_io_s),
    .io_cout(m_2339_io_cout)
  );
  Adder m_2340 ( // @[MUL.scala 102:19]
    .io_x1(m_2340_io_x1),
    .io_x2(m_2340_io_x2),
    .io_x3(m_2340_io_x3),
    .io_s(m_2340_io_s),
    .io_cout(m_2340_io_cout)
  );
  Adder m_2341 ( // @[MUL.scala 102:19]
    .io_x1(m_2341_io_x1),
    .io_x2(m_2341_io_x2),
    .io_x3(m_2341_io_x3),
    .io_s(m_2341_io_s),
    .io_cout(m_2341_io_cout)
  );
  Adder m_2342 ( // @[MUL.scala 102:19]
    .io_x1(m_2342_io_x1),
    .io_x2(m_2342_io_x2),
    .io_x3(m_2342_io_x3),
    .io_s(m_2342_io_s),
    .io_cout(m_2342_io_cout)
  );
  Adder m_2343 ( // @[MUL.scala 102:19]
    .io_x1(m_2343_io_x1),
    .io_x2(m_2343_io_x2),
    .io_x3(m_2343_io_x3),
    .io_s(m_2343_io_s),
    .io_cout(m_2343_io_cout)
  );
  Adder m_2344 ( // @[MUL.scala 102:19]
    .io_x1(m_2344_io_x1),
    .io_x2(m_2344_io_x2),
    .io_x3(m_2344_io_x3),
    .io_s(m_2344_io_s),
    .io_cout(m_2344_io_cout)
  );
  Adder m_2345 ( // @[MUL.scala 102:19]
    .io_x1(m_2345_io_x1),
    .io_x2(m_2345_io_x2),
    .io_x3(m_2345_io_x3),
    .io_s(m_2345_io_s),
    .io_cout(m_2345_io_cout)
  );
  Adder m_2346 ( // @[MUL.scala 102:19]
    .io_x1(m_2346_io_x1),
    .io_x2(m_2346_io_x2),
    .io_x3(m_2346_io_x3),
    .io_s(m_2346_io_s),
    .io_cout(m_2346_io_cout)
  );
  Adder m_2347 ( // @[MUL.scala 102:19]
    .io_x1(m_2347_io_x1),
    .io_x2(m_2347_io_x2),
    .io_x3(m_2347_io_x3),
    .io_s(m_2347_io_s),
    .io_cout(m_2347_io_cout)
  );
  Adder m_2348 ( // @[MUL.scala 102:19]
    .io_x1(m_2348_io_x1),
    .io_x2(m_2348_io_x2),
    .io_x3(m_2348_io_x3),
    .io_s(m_2348_io_s),
    .io_cout(m_2348_io_cout)
  );
  Adder m_2349 ( // @[MUL.scala 102:19]
    .io_x1(m_2349_io_x1),
    .io_x2(m_2349_io_x2),
    .io_x3(m_2349_io_x3),
    .io_s(m_2349_io_s),
    .io_cout(m_2349_io_cout)
  );
  Adder m_2350 ( // @[MUL.scala 102:19]
    .io_x1(m_2350_io_x1),
    .io_x2(m_2350_io_x2),
    .io_x3(m_2350_io_x3),
    .io_s(m_2350_io_s),
    .io_cout(m_2350_io_cout)
  );
  Adder m_2351 ( // @[MUL.scala 102:19]
    .io_x1(m_2351_io_x1),
    .io_x2(m_2351_io_x2),
    .io_x3(m_2351_io_x3),
    .io_s(m_2351_io_s),
    .io_cout(m_2351_io_cout)
  );
  Adder m_2352 ( // @[MUL.scala 102:19]
    .io_x1(m_2352_io_x1),
    .io_x2(m_2352_io_x2),
    .io_x3(m_2352_io_x3),
    .io_s(m_2352_io_s),
    .io_cout(m_2352_io_cout)
  );
  Adder m_2353 ( // @[MUL.scala 102:19]
    .io_x1(m_2353_io_x1),
    .io_x2(m_2353_io_x2),
    .io_x3(m_2353_io_x3),
    .io_s(m_2353_io_s),
    .io_cout(m_2353_io_cout)
  );
  Adder m_2354 ( // @[MUL.scala 102:19]
    .io_x1(m_2354_io_x1),
    .io_x2(m_2354_io_x2),
    .io_x3(m_2354_io_x3),
    .io_s(m_2354_io_s),
    .io_cout(m_2354_io_cout)
  );
  Adder m_2355 ( // @[MUL.scala 102:19]
    .io_x1(m_2355_io_x1),
    .io_x2(m_2355_io_x2),
    .io_x3(m_2355_io_x3),
    .io_s(m_2355_io_s),
    .io_cout(m_2355_io_cout)
  );
  Adder m_2356 ( // @[MUL.scala 102:19]
    .io_x1(m_2356_io_x1),
    .io_x2(m_2356_io_x2),
    .io_x3(m_2356_io_x3),
    .io_s(m_2356_io_s),
    .io_cout(m_2356_io_cout)
  );
  Adder m_2357 ( // @[MUL.scala 102:19]
    .io_x1(m_2357_io_x1),
    .io_x2(m_2357_io_x2),
    .io_x3(m_2357_io_x3),
    .io_s(m_2357_io_s),
    .io_cout(m_2357_io_cout)
  );
  Adder m_2358 ( // @[MUL.scala 102:19]
    .io_x1(m_2358_io_x1),
    .io_x2(m_2358_io_x2),
    .io_x3(m_2358_io_x3),
    .io_s(m_2358_io_s),
    .io_cout(m_2358_io_cout)
  );
  Adder m_2359 ( // @[MUL.scala 102:19]
    .io_x1(m_2359_io_x1),
    .io_x2(m_2359_io_x2),
    .io_x3(m_2359_io_x3),
    .io_s(m_2359_io_s),
    .io_cout(m_2359_io_cout)
  );
  Adder m_2360 ( // @[MUL.scala 102:19]
    .io_x1(m_2360_io_x1),
    .io_x2(m_2360_io_x2),
    .io_x3(m_2360_io_x3),
    .io_s(m_2360_io_s),
    .io_cout(m_2360_io_cout)
  );
  Adder m_2361 ( // @[MUL.scala 102:19]
    .io_x1(m_2361_io_x1),
    .io_x2(m_2361_io_x2),
    .io_x3(m_2361_io_x3),
    .io_s(m_2361_io_s),
    .io_cout(m_2361_io_cout)
  );
  Adder m_2362 ( // @[MUL.scala 102:19]
    .io_x1(m_2362_io_x1),
    .io_x2(m_2362_io_x2),
    .io_x3(m_2362_io_x3),
    .io_s(m_2362_io_s),
    .io_cout(m_2362_io_cout)
  );
  Adder m_2363 ( // @[MUL.scala 102:19]
    .io_x1(m_2363_io_x1),
    .io_x2(m_2363_io_x2),
    .io_x3(m_2363_io_x3),
    .io_s(m_2363_io_s),
    .io_cout(m_2363_io_cout)
  );
  Adder m_2364 ( // @[MUL.scala 102:19]
    .io_x1(m_2364_io_x1),
    .io_x2(m_2364_io_x2),
    .io_x3(m_2364_io_x3),
    .io_s(m_2364_io_s),
    .io_cout(m_2364_io_cout)
  );
  Adder m_2365 ( // @[MUL.scala 102:19]
    .io_x1(m_2365_io_x1),
    .io_x2(m_2365_io_x2),
    .io_x3(m_2365_io_x3),
    .io_s(m_2365_io_s),
    .io_cout(m_2365_io_cout)
  );
  Adder m_2366 ( // @[MUL.scala 102:19]
    .io_x1(m_2366_io_x1),
    .io_x2(m_2366_io_x2),
    .io_x3(m_2366_io_x3),
    .io_s(m_2366_io_s),
    .io_cout(m_2366_io_cout)
  );
  Adder m_2367 ( // @[MUL.scala 102:19]
    .io_x1(m_2367_io_x1),
    .io_x2(m_2367_io_x2),
    .io_x3(m_2367_io_x3),
    .io_s(m_2367_io_s),
    .io_cout(m_2367_io_cout)
  );
  Adder m_2368 ( // @[MUL.scala 102:19]
    .io_x1(m_2368_io_x1),
    .io_x2(m_2368_io_x2),
    .io_x3(m_2368_io_x3),
    .io_s(m_2368_io_s),
    .io_cout(m_2368_io_cout)
  );
  Adder m_2369 ( // @[MUL.scala 102:19]
    .io_x1(m_2369_io_x1),
    .io_x2(m_2369_io_x2),
    .io_x3(m_2369_io_x3),
    .io_s(m_2369_io_s),
    .io_cout(m_2369_io_cout)
  );
  Adder m_2370 ( // @[MUL.scala 102:19]
    .io_x1(m_2370_io_x1),
    .io_x2(m_2370_io_x2),
    .io_x3(m_2370_io_x3),
    .io_s(m_2370_io_s),
    .io_cout(m_2370_io_cout)
  );
  Adder m_2371 ( // @[MUL.scala 102:19]
    .io_x1(m_2371_io_x1),
    .io_x2(m_2371_io_x2),
    .io_x3(m_2371_io_x3),
    .io_s(m_2371_io_s),
    .io_cout(m_2371_io_cout)
  );
  Adder m_2372 ( // @[MUL.scala 102:19]
    .io_x1(m_2372_io_x1),
    .io_x2(m_2372_io_x2),
    .io_x3(m_2372_io_x3),
    .io_s(m_2372_io_s),
    .io_cout(m_2372_io_cout)
  );
  Adder m_2373 ( // @[MUL.scala 102:19]
    .io_x1(m_2373_io_x1),
    .io_x2(m_2373_io_x2),
    .io_x3(m_2373_io_x3),
    .io_s(m_2373_io_s),
    .io_cout(m_2373_io_cout)
  );
  Adder m_2374 ( // @[MUL.scala 102:19]
    .io_x1(m_2374_io_x1),
    .io_x2(m_2374_io_x2),
    .io_x3(m_2374_io_x3),
    .io_s(m_2374_io_s),
    .io_cout(m_2374_io_cout)
  );
  Adder m_2375 ( // @[MUL.scala 102:19]
    .io_x1(m_2375_io_x1),
    .io_x2(m_2375_io_x2),
    .io_x3(m_2375_io_x3),
    .io_s(m_2375_io_s),
    .io_cout(m_2375_io_cout)
  );
  Adder m_2376 ( // @[MUL.scala 102:19]
    .io_x1(m_2376_io_x1),
    .io_x2(m_2376_io_x2),
    .io_x3(m_2376_io_x3),
    .io_s(m_2376_io_s),
    .io_cout(m_2376_io_cout)
  );
  Half_Adder m_2377 ( // @[MUL.scala 124:19]
    .io_in_0(m_2377_io_in_0),
    .io_in_1(m_2377_io_in_1),
    .io_out_0(m_2377_io_out_0),
    .io_out_1(m_2377_io_out_1)
  );
  Half_Adder m_2378 ( // @[MUL.scala 124:19]
    .io_in_0(m_2378_io_in_0),
    .io_in_1(m_2378_io_in_1),
    .io_out_0(m_2378_io_out_0),
    .io_out_1(m_2378_io_out_1)
  );
  Half_Adder m_2379 ( // @[MUL.scala 124:19]
    .io_in_0(m_2379_io_in_0),
    .io_in_1(m_2379_io_in_1),
    .io_out_0(m_2379_io_out_0),
    .io_out_1(m_2379_io_out_1)
  );
  Half_Adder m_2380 ( // @[MUL.scala 124:19]
    .io_in_0(m_2380_io_in_0),
    .io_in_1(m_2380_io_in_1),
    .io_out_0(m_2380_io_out_0),
    .io_out_1(m_2380_io_out_1)
  );
  Half_Adder m_2381 ( // @[MUL.scala 124:19]
    .io_in_0(m_2381_io_in_0),
    .io_in_1(m_2381_io_in_1),
    .io_out_0(m_2381_io_out_0),
    .io_out_1(m_2381_io_out_1)
  );
  Half_Adder m_2382 ( // @[MUL.scala 124:19]
    .io_in_0(m_2382_io_in_0),
    .io_in_1(m_2382_io_in_1),
    .io_out_0(m_2382_io_out_0),
    .io_out_1(m_2382_io_out_1)
  );
  Half_Adder m_2383 ( // @[MUL.scala 124:19]
    .io_in_0(m_2383_io_in_0),
    .io_in_1(m_2383_io_in_1),
    .io_out_0(m_2383_io_out_0),
    .io_out_1(m_2383_io_out_1)
  );
  Half_Adder m_2384 ( // @[MUL.scala 124:19]
    .io_in_0(m_2384_io_in_0),
    .io_in_1(m_2384_io_in_1),
    .io_out_0(m_2384_io_out_0),
    .io_out_1(m_2384_io_out_1)
  );
  Half_Adder m_2385 ( // @[MUL.scala 124:19]
    .io_in_0(m_2385_io_in_0),
    .io_in_1(m_2385_io_in_1),
    .io_out_0(m_2385_io_out_0),
    .io_out_1(m_2385_io_out_1)
  );
  Half_Adder m_2386 ( // @[MUL.scala 124:19]
    .io_in_0(m_2386_io_in_0),
    .io_in_1(m_2386_io_in_1),
    .io_out_0(m_2386_io_out_0),
    .io_out_1(m_2386_io_out_1)
  );
  Half_Adder m_2387 ( // @[MUL.scala 124:19]
    .io_in_0(m_2387_io_in_0),
    .io_in_1(m_2387_io_in_1),
    .io_out_0(m_2387_io_out_0),
    .io_out_1(m_2387_io_out_1)
  );
  Half_Adder m_2388 ( // @[MUL.scala 124:19]
    .io_in_0(m_2388_io_in_0),
    .io_in_1(m_2388_io_in_1),
    .io_out_0(m_2388_io_out_0),
    .io_out_1(m_2388_io_out_1)
  );
  Half_Adder m_2389 ( // @[MUL.scala 124:19]
    .io_in_0(m_2389_io_in_0),
    .io_in_1(m_2389_io_in_1),
    .io_out_0(m_2389_io_out_0),
    .io_out_1(m_2389_io_out_1)
  );
  Half_Adder m_2390 ( // @[MUL.scala 124:19]
    .io_in_0(m_2390_io_in_0),
    .io_in_1(m_2390_io_in_1),
    .io_out_0(m_2390_io_out_0),
    .io_out_1(m_2390_io_out_1)
  );
  Half_Adder m_2391 ( // @[MUL.scala 124:19]
    .io_in_0(m_2391_io_in_0),
    .io_in_1(m_2391_io_in_1),
    .io_out_0(m_2391_io_out_0),
    .io_out_1(m_2391_io_out_1)
  );
  Half_Adder m_2392 ( // @[MUL.scala 124:19]
    .io_in_0(m_2392_io_in_0),
    .io_in_1(m_2392_io_in_1),
    .io_out_0(m_2392_io_out_0),
    .io_out_1(m_2392_io_out_1)
  );
  Half_Adder m_2393 ( // @[MUL.scala 124:19]
    .io_in_0(m_2393_io_in_0),
    .io_in_1(m_2393_io_in_1),
    .io_out_0(m_2393_io_out_0),
    .io_out_1(m_2393_io_out_1)
  );
  Half_Adder m_2394 ( // @[MUL.scala 124:19]
    .io_in_0(m_2394_io_in_0),
    .io_in_1(m_2394_io_in_1),
    .io_out_0(m_2394_io_out_0),
    .io_out_1(m_2394_io_out_1)
  );
  Half_Adder m_2395 ( // @[MUL.scala 124:19]
    .io_in_0(m_2395_io_in_0),
    .io_in_1(m_2395_io_in_1),
    .io_out_0(m_2395_io_out_0),
    .io_out_1(m_2395_io_out_1)
  );
  Half_Adder m_2396 ( // @[MUL.scala 124:19]
    .io_in_0(m_2396_io_in_0),
    .io_in_1(m_2396_io_in_1),
    .io_out_0(m_2396_io_out_0),
    .io_out_1(m_2396_io_out_1)
  );
  Half_Adder m_2397 ( // @[MUL.scala 124:19]
    .io_in_0(m_2397_io_in_0),
    .io_in_1(m_2397_io_in_1),
    .io_out_0(m_2397_io_out_0),
    .io_out_1(m_2397_io_out_1)
  );
  Half_Adder m_2398 ( // @[MUL.scala 124:19]
    .io_in_0(m_2398_io_in_0),
    .io_in_1(m_2398_io_in_1),
    .io_out_0(m_2398_io_out_0),
    .io_out_1(m_2398_io_out_1)
  );
  Half_Adder m_2399 ( // @[MUL.scala 124:19]
    .io_in_0(m_2399_io_in_0),
    .io_in_1(m_2399_io_in_1),
    .io_out_0(m_2399_io_out_0),
    .io_out_1(m_2399_io_out_1)
  );
  Half_Adder m_2400 ( // @[MUL.scala 124:19]
    .io_in_0(m_2400_io_in_0),
    .io_in_1(m_2400_io_in_1),
    .io_out_0(m_2400_io_out_0),
    .io_out_1(m_2400_io_out_1)
  );
  Half_Adder m_2401 ( // @[MUL.scala 124:19]
    .io_in_0(m_2401_io_in_0),
    .io_in_1(m_2401_io_in_1),
    .io_out_0(m_2401_io_out_0),
    .io_out_1(m_2401_io_out_1)
  );
  Half_Adder m_2402 ( // @[MUL.scala 124:19]
    .io_in_0(m_2402_io_in_0),
    .io_in_1(m_2402_io_in_1),
    .io_out_0(m_2402_io_out_0),
    .io_out_1(m_2402_io_out_1)
  );
  Half_Adder m_2403 ( // @[MUL.scala 124:19]
    .io_in_0(m_2403_io_in_0),
    .io_in_1(m_2403_io_in_1),
    .io_out_0(m_2403_io_out_0),
    .io_out_1(m_2403_io_out_1)
  );
  Half_Adder m_2404 ( // @[MUL.scala 124:19]
    .io_in_0(m_2404_io_in_0),
    .io_in_1(m_2404_io_in_1),
    .io_out_0(m_2404_io_out_0),
    .io_out_1(m_2404_io_out_1)
  );
  Half_Adder m_2405 ( // @[MUL.scala 124:19]
    .io_in_0(m_2405_io_in_0),
    .io_in_1(m_2405_io_in_1),
    .io_out_0(m_2405_io_out_0),
    .io_out_1(m_2405_io_out_1)
  );
  Half_Adder m_2406 ( // @[MUL.scala 124:19]
    .io_in_0(m_2406_io_in_0),
    .io_in_1(m_2406_io_in_1),
    .io_out_0(m_2406_io_out_0),
    .io_out_1(m_2406_io_out_1)
  );
  Half_Adder m_2407 ( // @[MUL.scala 124:19]
    .io_in_0(m_2407_io_in_0),
    .io_in_1(m_2407_io_in_1),
    .io_out_0(m_2407_io_out_0),
    .io_out_1(m_2407_io_out_1)
  );
  Half_Adder m_2408 ( // @[MUL.scala 124:19]
    .io_in_0(m_2408_io_in_0),
    .io_in_1(m_2408_io_in_1),
    .io_out_0(m_2408_io_out_0),
    .io_out_1(m_2408_io_out_1)
  );
  Half_Adder m_2409 ( // @[MUL.scala 124:19]
    .io_in_0(m_2409_io_in_0),
    .io_in_1(m_2409_io_in_1),
    .io_out_0(m_2409_io_out_0),
    .io_out_1(m_2409_io_out_1)
  );
  Half_Adder m_2410 ( // @[MUL.scala 124:19]
    .io_in_0(m_2410_io_in_0),
    .io_in_1(m_2410_io_in_1),
    .io_out_0(m_2410_io_out_0),
    .io_out_1(m_2410_io_out_1)
  );
  Half_Adder m_2411 ( // @[MUL.scala 124:19]
    .io_in_0(m_2411_io_in_0),
    .io_in_1(m_2411_io_in_1),
    .io_out_0(m_2411_io_out_0),
    .io_out_1(m_2411_io_out_1)
  );
  Half_Adder m_2412 ( // @[MUL.scala 124:19]
    .io_in_0(m_2412_io_in_0),
    .io_in_1(m_2412_io_in_1),
    .io_out_0(m_2412_io_out_0),
    .io_out_1(m_2412_io_out_1)
  );
  Half_Adder m_2413 ( // @[MUL.scala 124:19]
    .io_in_0(m_2413_io_in_0),
    .io_in_1(m_2413_io_in_1),
    .io_out_0(m_2413_io_out_0),
    .io_out_1(m_2413_io_out_1)
  );
  Half_Adder m_2414 ( // @[MUL.scala 124:19]
    .io_in_0(m_2414_io_in_0),
    .io_in_1(m_2414_io_in_1),
    .io_out_0(m_2414_io_out_0),
    .io_out_1(m_2414_io_out_1)
  );
  Half_Adder m_2415 ( // @[MUL.scala 124:19]
    .io_in_0(m_2415_io_in_0),
    .io_in_1(m_2415_io_in_1),
    .io_out_0(m_2415_io_out_0),
    .io_out_1(m_2415_io_out_1)
  );
  Half_Adder m_2416 ( // @[MUL.scala 124:19]
    .io_in_0(m_2416_io_in_0),
    .io_in_1(m_2416_io_in_1),
    .io_out_0(m_2416_io_out_0),
    .io_out_1(m_2416_io_out_1)
  );
  Half_Adder m_2417 ( // @[MUL.scala 124:19]
    .io_in_0(m_2417_io_in_0),
    .io_in_1(m_2417_io_in_1),
    .io_out_0(m_2417_io_out_0),
    .io_out_1(m_2417_io_out_1)
  );
  Half_Adder m_2418 ( // @[MUL.scala 124:19]
    .io_in_0(m_2418_io_in_0),
    .io_in_1(m_2418_io_in_1),
    .io_out_0(m_2418_io_out_0),
    .io_out_1(m_2418_io_out_1)
  );
  Half_Adder m_2419 ( // @[MUL.scala 124:19]
    .io_in_0(m_2419_io_in_0),
    .io_in_1(m_2419_io_in_1),
    .io_out_0(m_2419_io_out_0),
    .io_out_1(m_2419_io_out_1)
  );
  Half_Adder m_2420 ( // @[MUL.scala 124:19]
    .io_in_0(m_2420_io_in_0),
    .io_in_1(m_2420_io_in_1),
    .io_out_0(m_2420_io_out_0),
    .io_out_1(m_2420_io_out_1)
  );
  Half_Adder m_2421 ( // @[MUL.scala 124:19]
    .io_in_0(m_2421_io_in_0),
    .io_in_1(m_2421_io_in_1),
    .io_out_0(m_2421_io_out_0),
    .io_out_1(m_2421_io_out_1)
  );
  Half_Adder m_2422 ( // @[MUL.scala 124:19]
    .io_in_0(m_2422_io_in_0),
    .io_in_1(m_2422_io_in_1),
    .io_out_0(m_2422_io_out_0),
    .io_out_1(m_2422_io_out_1)
  );
  Half_Adder m_2423 ( // @[MUL.scala 124:19]
    .io_in_0(m_2423_io_in_0),
    .io_in_1(m_2423_io_in_1),
    .io_out_0(m_2423_io_out_0),
    .io_out_1(m_2423_io_out_1)
  );
  Half_Adder m_2424 ( // @[MUL.scala 124:19]
    .io_in_0(m_2424_io_in_0),
    .io_in_1(m_2424_io_in_1),
    .io_out_0(m_2424_io_out_0),
    .io_out_1(m_2424_io_out_1)
  );
  Half_Adder m_2425 ( // @[MUL.scala 124:19]
    .io_in_0(m_2425_io_in_0),
    .io_in_1(m_2425_io_in_1),
    .io_out_0(m_2425_io_out_0),
    .io_out_1(m_2425_io_out_1)
  );
  Half_Adder m_2426 ( // @[MUL.scala 124:19]
    .io_in_0(m_2426_io_in_0),
    .io_in_1(m_2426_io_in_1),
    .io_out_0(m_2426_io_out_0),
    .io_out_1(m_2426_io_out_1)
  );
  Half_Adder m_2427 ( // @[MUL.scala 124:19]
    .io_in_0(m_2427_io_in_0),
    .io_in_1(m_2427_io_in_1),
    .io_out_0(m_2427_io_out_0),
    .io_out_1(m_2427_io_out_1)
  );
  Half_Adder m_2428 ( // @[MUL.scala 124:19]
    .io_in_0(m_2428_io_in_0),
    .io_in_1(m_2428_io_in_1),
    .io_out_0(m_2428_io_out_0),
    .io_out_1(m_2428_io_out_1)
  );
  Half_Adder m_2429 ( // @[MUL.scala 124:19]
    .io_in_0(m_2429_io_in_0),
    .io_in_1(m_2429_io_in_1),
    .io_out_0(m_2429_io_out_0),
    .io_out_1(m_2429_io_out_1)
  );
  Half_Adder m_2430 ( // @[MUL.scala 124:19]
    .io_in_0(m_2430_io_in_0),
    .io_in_1(m_2430_io_in_1),
    .io_out_0(m_2430_io_out_0),
    .io_out_1(m_2430_io_out_1)
  );
  Half_Adder m_2431 ( // @[MUL.scala 124:19]
    .io_in_0(m_2431_io_in_0),
    .io_in_1(m_2431_io_in_1),
    .io_out_0(m_2431_io_out_0),
    .io_out_1(m_2431_io_out_1)
  );
  Half_Adder m_2432 ( // @[MUL.scala 124:19]
    .io_in_0(m_2432_io_in_0),
    .io_in_1(m_2432_io_in_1),
    .io_out_0(m_2432_io_out_0),
    .io_out_1(m_2432_io_out_1)
  );
  Half_Adder m_2433 ( // @[MUL.scala 124:19]
    .io_in_0(m_2433_io_in_0),
    .io_in_1(m_2433_io_in_1),
    .io_out_0(m_2433_io_out_0),
    .io_out_1(m_2433_io_out_1)
  );
  Half_Adder m_2434 ( // @[MUL.scala 124:19]
    .io_in_0(m_2434_io_in_0),
    .io_in_1(m_2434_io_in_1),
    .io_out_0(m_2434_io_out_0),
    .io_out_1(m_2434_io_out_1)
  );
  Half_Adder m_2435 ( // @[MUL.scala 124:19]
    .io_in_0(m_2435_io_in_0),
    .io_in_1(m_2435_io_in_1),
    .io_out_0(m_2435_io_out_0),
    .io_out_1(m_2435_io_out_1)
  );
  Half_Adder m_2436 ( // @[MUL.scala 124:19]
    .io_in_0(m_2436_io_in_0),
    .io_in_1(m_2436_io_in_1),
    .io_out_0(m_2436_io_out_0),
    .io_out_1(m_2436_io_out_1)
  );
  Half_Adder m_2437 ( // @[MUL.scala 124:19]
    .io_in_0(m_2437_io_in_0),
    .io_in_1(m_2437_io_in_1),
    .io_out_0(m_2437_io_out_0),
    .io_out_1(m_2437_io_out_1)
  );
  Half_Adder m_2438 ( // @[MUL.scala 124:19]
    .io_in_0(m_2438_io_in_0),
    .io_in_1(m_2438_io_in_1),
    .io_out_0(m_2438_io_out_0),
    .io_out_1(m_2438_io_out_1)
  );
  Half_Adder m_2439 ( // @[MUL.scala 124:19]
    .io_in_0(m_2439_io_in_0),
    .io_in_1(m_2439_io_in_1),
    .io_out_0(m_2439_io_out_0),
    .io_out_1(m_2439_io_out_1)
  );
  Half_Adder m_2440 ( // @[MUL.scala 124:19]
    .io_in_0(m_2440_io_in_0),
    .io_in_1(m_2440_io_in_1),
    .io_out_0(m_2440_io_out_0),
    .io_out_1(m_2440_io_out_1)
  );
  Half_Adder m_2441 ( // @[MUL.scala 124:19]
    .io_in_0(m_2441_io_in_0),
    .io_in_1(m_2441_io_in_1),
    .io_out_0(m_2441_io_out_0),
    .io_out_1(m_2441_io_out_1)
  );
  Half_Adder m_2442 ( // @[MUL.scala 124:19]
    .io_in_0(m_2442_io_in_0),
    .io_in_1(m_2442_io_in_1),
    .io_out_0(m_2442_io_out_0),
    .io_out_1(m_2442_io_out_1)
  );
  Half_Adder m_2443 ( // @[MUL.scala 124:19]
    .io_in_0(m_2443_io_in_0),
    .io_in_1(m_2443_io_in_1),
    .io_out_0(m_2443_io_out_0),
    .io_out_1(m_2443_io_out_1)
  );
  Half_Adder m_2444 ( // @[MUL.scala 124:19]
    .io_in_0(m_2444_io_in_0),
    .io_in_1(m_2444_io_in_1),
    .io_out_0(m_2444_io_out_0),
    .io_out_1(m_2444_io_out_1)
  );
  Half_Adder m_2445 ( // @[MUL.scala 124:19]
    .io_in_0(m_2445_io_in_0),
    .io_in_1(m_2445_io_in_1),
    .io_out_0(m_2445_io_out_0),
    .io_out_1(m_2445_io_out_1)
  );
  Half_Adder m_2446 ( // @[MUL.scala 124:19]
    .io_in_0(m_2446_io_in_0),
    .io_in_1(m_2446_io_in_1),
    .io_out_0(m_2446_io_out_0),
    .io_out_1(m_2446_io_out_1)
  );
  Half_Adder m_2447 ( // @[MUL.scala 124:19]
    .io_in_0(m_2447_io_in_0),
    .io_in_1(m_2447_io_in_1),
    .io_out_0(m_2447_io_out_0),
    .io_out_1(m_2447_io_out_1)
  );
  Half_Adder m_2448 ( // @[MUL.scala 124:19]
    .io_in_0(m_2448_io_in_0),
    .io_in_1(m_2448_io_in_1),
    .io_out_0(m_2448_io_out_0),
    .io_out_1(m_2448_io_out_1)
  );
  Half_Adder m_2449 ( // @[MUL.scala 124:19]
    .io_in_0(m_2449_io_in_0),
    .io_in_1(m_2449_io_in_1),
    .io_out_0(m_2449_io_out_0),
    .io_out_1(m_2449_io_out_1)
  );
  Half_Adder m_2450 ( // @[MUL.scala 124:19]
    .io_in_0(m_2450_io_in_0),
    .io_in_1(m_2450_io_in_1),
    .io_out_0(m_2450_io_out_0),
    .io_out_1(m_2450_io_out_1)
  );
  Half_Adder m_2451 ( // @[MUL.scala 124:19]
    .io_in_0(m_2451_io_in_0),
    .io_in_1(m_2451_io_in_1),
    .io_out_0(m_2451_io_out_0),
    .io_out_1(m_2451_io_out_1)
  );
  Half_Adder m_2452 ( // @[MUL.scala 124:19]
    .io_in_0(m_2452_io_in_0),
    .io_in_1(m_2452_io_in_1),
    .io_out_0(m_2452_io_out_0),
    .io_out_1(m_2452_io_out_1)
  );
  Half_Adder m_2453 ( // @[MUL.scala 124:19]
    .io_in_0(m_2453_io_in_0),
    .io_in_1(m_2453_io_in_1),
    .io_out_0(m_2453_io_out_0),
    .io_out_1(m_2453_io_out_1)
  );
  Half_Adder m_2454 ( // @[MUL.scala 124:19]
    .io_in_0(m_2454_io_in_0),
    .io_in_1(m_2454_io_in_1),
    .io_out_0(m_2454_io_out_0),
    .io_out_1(m_2454_io_out_1)
  );
  Half_Adder m_2455 ( // @[MUL.scala 124:19]
    .io_in_0(m_2455_io_in_0),
    .io_in_1(m_2455_io_in_1),
    .io_out_0(m_2455_io_out_0),
    .io_out_1(m_2455_io_out_1)
  );
  Half_Adder m_2456 ( // @[MUL.scala 124:19]
    .io_in_0(m_2456_io_in_0),
    .io_in_1(m_2456_io_in_1),
    .io_out_0(m_2456_io_out_0),
    .io_out_1(m_2456_io_out_1)
  );
  Half_Adder m_2457 ( // @[MUL.scala 124:19]
    .io_in_0(m_2457_io_in_0),
    .io_in_1(m_2457_io_in_1),
    .io_out_0(m_2457_io_out_0),
    .io_out_1(m_2457_io_out_1)
  );
  Half_Adder m_2458 ( // @[MUL.scala 124:19]
    .io_in_0(m_2458_io_in_0),
    .io_in_1(m_2458_io_in_1),
    .io_out_0(m_2458_io_out_0),
    .io_out_1(m_2458_io_out_1)
  );
  Half_Adder m_2459 ( // @[MUL.scala 124:19]
    .io_in_0(m_2459_io_in_0),
    .io_in_1(m_2459_io_in_1),
    .io_out_0(m_2459_io_out_0),
    .io_out_1(m_2459_io_out_1)
  );
  Half_Adder m_2460 ( // @[MUL.scala 124:19]
    .io_in_0(m_2460_io_in_0),
    .io_in_1(m_2460_io_in_1),
    .io_out_0(m_2460_io_out_0),
    .io_out_1(m_2460_io_out_1)
  );
  Half_Adder m_2461 ( // @[MUL.scala 124:19]
    .io_in_0(m_2461_io_in_0),
    .io_in_1(m_2461_io_in_1),
    .io_out_0(m_2461_io_out_0),
    .io_out_1(m_2461_io_out_1)
  );
  Adder m_2462 ( // @[MUL.scala 102:19]
    .io_x1(m_2462_io_x1),
    .io_x2(m_2462_io_x2),
    .io_x3(m_2462_io_x3),
    .io_s(m_2462_io_s),
    .io_cout(m_2462_io_cout)
  );
  Adder m_2463 ( // @[MUL.scala 102:19]
    .io_x1(m_2463_io_x1),
    .io_x2(m_2463_io_x2),
    .io_x3(m_2463_io_x3),
    .io_s(m_2463_io_s),
    .io_cout(m_2463_io_cout)
  );
  Adder m_2464 ( // @[MUL.scala 102:19]
    .io_x1(m_2464_io_x1),
    .io_x2(m_2464_io_x2),
    .io_x3(m_2464_io_x3),
    .io_s(m_2464_io_s),
    .io_cout(m_2464_io_cout)
  );
  Adder m_2465 ( // @[MUL.scala 102:19]
    .io_x1(m_2465_io_x1),
    .io_x2(m_2465_io_x2),
    .io_x3(m_2465_io_x3),
    .io_s(m_2465_io_s),
    .io_cout(m_2465_io_cout)
  );
  Adder m_2466 ( // @[MUL.scala 102:19]
    .io_x1(m_2466_io_x1),
    .io_x2(m_2466_io_x2),
    .io_x3(m_2466_io_x3),
    .io_s(m_2466_io_s),
    .io_cout(m_2466_io_cout)
  );
  Adder m_2467 ( // @[MUL.scala 102:19]
    .io_x1(m_2467_io_x1),
    .io_x2(m_2467_io_x2),
    .io_x3(m_2467_io_x3),
    .io_s(m_2467_io_s),
    .io_cout(m_2467_io_cout)
  );
  Adder m_2468 ( // @[MUL.scala 102:19]
    .io_x1(m_2468_io_x1),
    .io_x2(m_2468_io_x2),
    .io_x3(m_2468_io_x3),
    .io_s(m_2468_io_s),
    .io_cout(m_2468_io_cout)
  );
  Adder m_2469 ( // @[MUL.scala 102:19]
    .io_x1(m_2469_io_x1),
    .io_x2(m_2469_io_x2),
    .io_x3(m_2469_io_x3),
    .io_s(m_2469_io_s),
    .io_cout(m_2469_io_cout)
  );
  Adder m_2470 ( // @[MUL.scala 102:19]
    .io_x1(m_2470_io_x1),
    .io_x2(m_2470_io_x2),
    .io_x3(m_2470_io_x3),
    .io_s(m_2470_io_s),
    .io_cout(m_2470_io_cout)
  );
  Adder m_2471 ( // @[MUL.scala 102:19]
    .io_x1(m_2471_io_x1),
    .io_x2(m_2471_io_x2),
    .io_x3(m_2471_io_x3),
    .io_s(m_2471_io_s),
    .io_cout(m_2471_io_cout)
  );
  Adder m_2472 ( // @[MUL.scala 102:19]
    .io_x1(m_2472_io_x1),
    .io_x2(m_2472_io_x2),
    .io_x3(m_2472_io_x3),
    .io_s(m_2472_io_s),
    .io_cout(m_2472_io_cout)
  );
  Adder m_2473 ( // @[MUL.scala 102:19]
    .io_x1(m_2473_io_x1),
    .io_x2(m_2473_io_x2),
    .io_x3(m_2473_io_x3),
    .io_s(m_2473_io_s),
    .io_cout(m_2473_io_cout)
  );
  Adder m_2474 ( // @[MUL.scala 102:19]
    .io_x1(m_2474_io_x1),
    .io_x2(m_2474_io_x2),
    .io_x3(m_2474_io_x3),
    .io_s(m_2474_io_s),
    .io_cout(m_2474_io_cout)
  );
  Adder m_2475 ( // @[MUL.scala 102:19]
    .io_x1(m_2475_io_x1),
    .io_x2(m_2475_io_x2),
    .io_x3(m_2475_io_x3),
    .io_s(m_2475_io_s),
    .io_cout(m_2475_io_cout)
  );
  Adder m_2476 ( // @[MUL.scala 102:19]
    .io_x1(m_2476_io_x1),
    .io_x2(m_2476_io_x2),
    .io_x3(m_2476_io_x3),
    .io_s(m_2476_io_s),
    .io_cout(m_2476_io_cout)
  );
  Adder m_2477 ( // @[MUL.scala 102:19]
    .io_x1(m_2477_io_x1),
    .io_x2(m_2477_io_x2),
    .io_x3(m_2477_io_x3),
    .io_s(m_2477_io_s),
    .io_cout(m_2477_io_cout)
  );
  Adder m_2478 ( // @[MUL.scala 102:19]
    .io_x1(m_2478_io_x1),
    .io_x2(m_2478_io_x2),
    .io_x3(m_2478_io_x3),
    .io_s(m_2478_io_s),
    .io_cout(m_2478_io_cout)
  );
  Adder m_2479 ( // @[MUL.scala 102:19]
    .io_x1(m_2479_io_x1),
    .io_x2(m_2479_io_x2),
    .io_x3(m_2479_io_x3),
    .io_s(m_2479_io_s),
    .io_cout(m_2479_io_cout)
  );
  Adder m_2480 ( // @[MUL.scala 102:19]
    .io_x1(m_2480_io_x1),
    .io_x2(m_2480_io_x2),
    .io_x3(m_2480_io_x3),
    .io_s(m_2480_io_s),
    .io_cout(m_2480_io_cout)
  );
  Adder m_2481 ( // @[MUL.scala 102:19]
    .io_x1(m_2481_io_x1),
    .io_x2(m_2481_io_x2),
    .io_x3(m_2481_io_x3),
    .io_s(m_2481_io_s),
    .io_cout(m_2481_io_cout)
  );
  Adder m_2482 ( // @[MUL.scala 102:19]
    .io_x1(m_2482_io_x1),
    .io_x2(m_2482_io_x2),
    .io_x3(m_2482_io_x3),
    .io_s(m_2482_io_s),
    .io_cout(m_2482_io_cout)
  );
  Half_Adder m_2483 ( // @[MUL.scala 124:19]
    .io_in_0(m_2483_io_in_0),
    .io_in_1(m_2483_io_in_1),
    .io_out_0(m_2483_io_out_0),
    .io_out_1(m_2483_io_out_1)
  );
  Half_Adder m_2484 ( // @[MUL.scala 124:19]
    .io_in_0(m_2484_io_in_0),
    .io_in_1(m_2484_io_in_1),
    .io_out_0(m_2484_io_out_0),
    .io_out_1(m_2484_io_out_1)
  );
  Half_Adder m_2485 ( // @[MUL.scala 124:19]
    .io_in_0(m_2485_io_in_0),
    .io_in_1(m_2485_io_in_1),
    .io_out_0(m_2485_io_out_0),
    .io_out_1(m_2485_io_out_1)
  );
  Half_Adder m_2486 ( // @[MUL.scala 124:19]
    .io_in_0(m_2486_io_in_0),
    .io_in_1(m_2486_io_in_1),
    .io_out_0(m_2486_io_out_0),
    .io_out_1(m_2486_io_out_1)
  );
  Half_Adder m_2487 ( // @[MUL.scala 124:19]
    .io_in_0(m_2487_io_in_0),
    .io_in_1(m_2487_io_in_1),
    .io_out_0(m_2487_io_out_0),
    .io_out_1(m_2487_io_out_1)
  );
  Half_Adder m_2488 ( // @[MUL.scala 124:19]
    .io_in_0(m_2488_io_in_0),
    .io_in_1(m_2488_io_in_1),
    .io_out_0(m_2488_io_out_0),
    .io_out_1(m_2488_io_out_1)
  );
  Half_Adder m_2489 ( // @[MUL.scala 124:19]
    .io_in_0(m_2489_io_in_0),
    .io_in_1(m_2489_io_in_1),
    .io_out_0(m_2489_io_out_0),
    .io_out_1(m_2489_io_out_1)
  );
  Half_Adder m_2490 ( // @[MUL.scala 124:19]
    .io_in_0(m_2490_io_in_0),
    .io_in_1(m_2490_io_in_1),
    .io_out_0(m_2490_io_out_0),
    .io_out_1(m_2490_io_out_1)
  );
  Half_Adder m_2491 ( // @[MUL.scala 124:19]
    .io_in_0(m_2491_io_in_0),
    .io_in_1(m_2491_io_in_1),
    .io_out_0(m_2491_io_out_0),
    .io_out_1(m_2491_io_out_1)
  );
  Half_Adder m_2492 ( // @[MUL.scala 124:19]
    .io_in_0(m_2492_io_in_0),
    .io_in_1(m_2492_io_in_1),
    .io_out_0(m_2492_io_out_0),
    .io_out_1(m_2492_io_out_1)
  );
  Half_Adder m_2493 ( // @[MUL.scala 124:19]
    .io_in_0(m_2493_io_in_0),
    .io_in_1(m_2493_io_in_1),
    .io_out_0(m_2493_io_out_0),
    .io_out_1(m_2493_io_out_1)
  );
  Half_Adder m_2494 ( // @[MUL.scala 124:19]
    .io_in_0(m_2494_io_in_0),
    .io_in_1(m_2494_io_in_1),
    .io_out_0(m_2494_io_out_0),
    .io_out_1(m_2494_io_out_1)
  );
  Half_Adder m_2495 ( // @[MUL.scala 124:19]
    .io_in_0(m_2495_io_in_0),
    .io_in_1(m_2495_io_in_1),
    .io_out_0(m_2495_io_out_0),
    .io_out_1(m_2495_io_out_1)
  );
  Half_Adder m_2496 ( // @[MUL.scala 124:19]
    .io_in_0(m_2496_io_in_0),
    .io_in_1(m_2496_io_in_1),
    .io_out_0(m_2496_io_out_0),
    .io_out_1(m_2496_io_out_1)
  );
  Half_Adder m_2497 ( // @[MUL.scala 124:19]
    .io_in_0(m_2497_io_in_0),
    .io_in_1(m_2497_io_in_1),
    .io_out_0(m_2497_io_out_0),
    .io_out_1(m_2497_io_out_1)
  );
  Half_Adder m_2498 ( // @[MUL.scala 124:19]
    .io_in_0(m_2498_io_in_0),
    .io_in_1(m_2498_io_in_1),
    .io_out_0(m_2498_io_out_0),
    .io_out_1(m_2498_io_out_1)
  );
  Half_Adder m_2499 ( // @[MUL.scala 124:19]
    .io_in_0(m_2499_io_in_0),
    .io_in_1(m_2499_io_in_1),
    .io_out_0(m_2499_io_out_0),
    .io_out_1(m_2499_io_out_1)
  );
  Half_Adder m_2500 ( // @[MUL.scala 124:19]
    .io_in_0(m_2500_io_in_0),
    .io_in_1(m_2500_io_in_1),
    .io_out_0(m_2500_io_out_0),
    .io_out_1(m_2500_io_out_1)
  );
  Half_Adder m_2501 ( // @[MUL.scala 124:19]
    .io_in_0(m_2501_io_in_0),
    .io_in_1(m_2501_io_in_1),
    .io_out_0(m_2501_io_out_0),
    .io_out_1(m_2501_io_out_1)
  );
  Half_Adder m_2502 ( // @[MUL.scala 124:19]
    .io_in_0(m_2502_io_in_0),
    .io_in_1(m_2502_io_in_1),
    .io_out_0(m_2502_io_out_0),
    .io_out_1(m_2502_io_out_1)
  );
  Half_Adder m_2503 ( // @[MUL.scala 124:19]
    .io_in_0(m_2503_io_in_0),
    .io_in_1(m_2503_io_in_1),
    .io_out_0(m_2503_io_out_0),
    .io_out_1(m_2503_io_out_1)
  );
  Half_Adder m_2504 ( // @[MUL.scala 124:19]
    .io_in_0(m_2504_io_in_0),
    .io_in_1(m_2504_io_in_1),
    .io_out_0(m_2504_io_out_0),
    .io_out_1(m_2504_io_out_1)
  );
  Half_Adder m_2505 ( // @[MUL.scala 124:19]
    .io_in_0(m_2505_io_in_0),
    .io_in_1(m_2505_io_in_1),
    .io_out_0(m_2505_io_out_0),
    .io_out_1(m_2505_io_out_1)
  );
  Half_Adder m_2506 ( // @[MUL.scala 124:19]
    .io_in_0(m_2506_io_in_0),
    .io_in_1(m_2506_io_in_1),
    .io_out_0(m_2506_io_out_0),
    .io_out_1(m_2506_io_out_1)
  );
  Half_Adder m_2507 ( // @[MUL.scala 124:19]
    .io_in_0(m_2507_io_in_0),
    .io_in_1(m_2507_io_in_1),
    .io_out_0(m_2507_io_out_0),
    .io_out_1(m_2507_io_out_1)
  );
  Half_Adder m_2508 ( // @[MUL.scala 124:19]
    .io_in_0(m_2508_io_in_0),
    .io_in_1(m_2508_io_in_1),
    .io_out_0(m_2508_io_out_0),
    .io_out_1(m_2508_io_out_1)
  );
  Half_Adder m_2509 ( // @[MUL.scala 124:19]
    .io_in_0(m_2509_io_in_0),
    .io_in_1(m_2509_io_in_1),
    .io_out_0(m_2509_io_out_0),
    .io_out_1(m_2509_io_out_1)
  );
  Half_Adder m_2510 ( // @[MUL.scala 124:19]
    .io_in_0(m_2510_io_in_0),
    .io_in_1(m_2510_io_in_1),
    .io_out_0(m_2510_io_out_0),
    .io_out_1(m_2510_io_out_1)
  );
  Half_Adder m_2511 ( // @[MUL.scala 124:19]
    .io_in_0(m_2511_io_in_0),
    .io_in_1(m_2511_io_in_1),
    .io_out_0(m_2511_io_out_0),
    .io_out_1(m_2511_io_out_1)
  );
  Half_Adder m_2512 ( // @[MUL.scala 124:19]
    .io_in_0(m_2512_io_in_0),
    .io_in_1(m_2512_io_in_1),
    .io_out_0(m_2512_io_out_0),
    .io_out_1(m_2512_io_out_1)
  );
  Half_Adder m_2513 ( // @[MUL.scala 124:19]
    .io_in_0(m_2513_io_in_0),
    .io_in_1(m_2513_io_in_1),
    .io_out_0(m_2513_io_out_0),
    .io_out_1(m_2513_io_out_1)
  );
  Half_Adder m_2514 ( // @[MUL.scala 124:19]
    .io_in_0(m_2514_io_in_0),
    .io_in_1(m_2514_io_in_1),
    .io_out_0(m_2514_io_out_0),
    .io_out_1(m_2514_io_out_1)
  );
  Half_Adder m_2515 ( // @[MUL.scala 124:19]
    .io_in_0(m_2515_io_in_0),
    .io_in_1(m_2515_io_in_1),
    .io_out_0(m_2515_io_out_0),
    .io_out_1(m_2515_io_out_1)
  );
  Half_Adder m_2516 ( // @[MUL.scala 124:19]
    .io_in_0(m_2516_io_in_0),
    .io_in_1(m_2516_io_in_1),
    .io_out_0(m_2516_io_out_0),
    .io_out_1(m_2516_io_out_1)
  );
  Half_Adder m_2517 ( // @[MUL.scala 124:19]
    .io_in_0(m_2517_io_in_0),
    .io_in_1(m_2517_io_in_1),
    .io_out_0(m_2517_io_out_0),
    .io_out_1(m_2517_io_out_1)
  );
  Half_Adder m_2518 ( // @[MUL.scala 124:19]
    .io_in_0(m_2518_io_in_0),
    .io_in_1(m_2518_io_in_1),
    .io_out_0(m_2518_io_out_0),
    .io_out_1(m_2518_io_out_1)
  );
  Half_Adder m_2519 ( // @[MUL.scala 124:19]
    .io_in_0(m_2519_io_in_0),
    .io_in_1(m_2519_io_in_1),
    .io_out_0(m_2519_io_out_0),
    .io_out_1(m_2519_io_out_1)
  );
  Half_Adder m_2520 ( // @[MUL.scala 124:19]
    .io_in_0(m_2520_io_in_0),
    .io_in_1(m_2520_io_in_1),
    .io_out_0(m_2520_io_out_0),
    .io_out_1(m_2520_io_out_1)
  );
  Half_Adder m_2521 ( // @[MUL.scala 124:19]
    .io_in_0(m_2521_io_in_0),
    .io_in_1(m_2521_io_in_1),
    .io_out_0(m_2521_io_out_0),
    .io_out_1(m_2521_io_out_1)
  );
  Half_Adder m_2522 ( // @[MUL.scala 124:19]
    .io_in_0(m_2522_io_in_0),
    .io_in_1(m_2522_io_in_1),
    .io_out_0(m_2522_io_out_0),
    .io_out_1(m_2522_io_out_1)
  );
  Half_Adder m_2523 ( // @[MUL.scala 124:19]
    .io_in_0(m_2523_io_in_0),
    .io_in_1(m_2523_io_in_1),
    .io_out_0(m_2523_io_out_0),
    .io_out_1(m_2523_io_out_1)
  );
  Half_Adder m_2524 ( // @[MUL.scala 124:19]
    .io_in_0(m_2524_io_in_0),
    .io_in_1(m_2524_io_in_1),
    .io_out_0(m_2524_io_out_0),
    .io_out_1(m_2524_io_out_1)
  );
  Half_Adder m_2525 ( // @[MUL.scala 124:19]
    .io_in_0(m_2525_io_in_0),
    .io_in_1(m_2525_io_in_1),
    .io_out_0(m_2525_io_out_0),
    .io_out_1(m_2525_io_out_1)
  );
  Half_Adder m_2526 ( // @[MUL.scala 124:19]
    .io_in_0(m_2526_io_in_0),
    .io_in_1(m_2526_io_in_1),
    .io_out_0(m_2526_io_out_0),
    .io_out_1(m_2526_io_out_1)
  );
  Half_Adder m_2527 ( // @[MUL.scala 124:19]
    .io_in_0(m_2527_io_in_0),
    .io_in_1(m_2527_io_in_1),
    .io_out_0(m_2527_io_out_0),
    .io_out_1(m_2527_io_out_1)
  );
  Half_Adder m_2528 ( // @[MUL.scala 124:19]
    .io_in_0(m_2528_io_in_0),
    .io_in_1(m_2528_io_in_1),
    .io_out_0(m_2528_io_out_0),
    .io_out_1(m_2528_io_out_1)
  );
  Half_Adder m_2529 ( // @[MUL.scala 124:19]
    .io_in_0(m_2529_io_in_0),
    .io_in_1(m_2529_io_in_1),
    .io_out_0(m_2529_io_out_0),
    .io_out_1(m_2529_io_out_1)
  );
  Half_Adder m_2530 ( // @[MUL.scala 124:19]
    .io_in_0(m_2530_io_in_0),
    .io_in_1(m_2530_io_in_1),
    .io_out_0(m_2530_io_out_0),
    .io_out_1(m_2530_io_out_1)
  );
  Half_Adder m_2531 ( // @[MUL.scala 124:19]
    .io_in_0(m_2531_io_in_0),
    .io_in_1(m_2531_io_in_1),
    .io_out_0(m_2531_io_out_0),
    .io_out_1(m_2531_io_out_1)
  );
  Half_Adder m_2532 ( // @[MUL.scala 124:19]
    .io_in_0(m_2532_io_in_0),
    .io_in_1(m_2532_io_in_1),
    .io_out_0(m_2532_io_out_0),
    .io_out_1(m_2532_io_out_1)
  );
  Half_Adder m_2533 ( // @[MUL.scala 124:19]
    .io_in_0(m_2533_io_in_0),
    .io_in_1(m_2533_io_in_1),
    .io_out_0(m_2533_io_out_0),
    .io_out_1(m_2533_io_out_1)
  );
  Half_Adder m_2534 ( // @[MUL.scala 124:19]
    .io_in_0(m_2534_io_in_0),
    .io_in_1(m_2534_io_in_1),
    .io_out_0(m_2534_io_out_0),
    .io_out_1(m_2534_io_out_1)
  );
  assign io_out_valid = count == 8'h2; // @[MUL.scala 335:17]
  assign io_out_bits_result_result_lo = result[63:0]; // @[MUL.scala 339:40]
  assign m_io_y_3 = src1[2:0]; // @[MUL.scala 303:56]
  assign m_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_1_io_y_3 = src1[4:2]; // @[MUL.scala 303:56]
  assign m_1_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_2_io_y_3 = src1[6:4]; // @[MUL.scala 303:56]
  assign m_2_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_3_io_y_3 = src1[8:6]; // @[MUL.scala 303:56]
  assign m_3_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_4_io_y_3 = src1[10:8]; // @[MUL.scala 303:56]
  assign m_4_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_5_io_y_3 = src1[12:10]; // @[MUL.scala 303:56]
  assign m_5_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_6_io_y_3 = src1[14:12]; // @[MUL.scala 303:56]
  assign m_6_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_7_io_y_3 = src1[16:14]; // @[MUL.scala 303:56]
  assign m_7_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_8_io_y_3 = src1[18:16]; // @[MUL.scala 303:56]
  assign m_8_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_9_io_y_3 = src1[20:18]; // @[MUL.scala 303:56]
  assign m_9_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_10_io_y_3 = src1[22:20]; // @[MUL.scala 303:56]
  assign m_10_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_11_io_y_3 = src1[24:22]; // @[MUL.scala 303:56]
  assign m_11_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_12_io_y_3 = src1[26:24]; // @[MUL.scala 303:56]
  assign m_12_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_13_io_y_3 = src1[28:26]; // @[MUL.scala 303:56]
  assign m_13_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_14_io_y_3 = src1[30:28]; // @[MUL.scala 303:56]
  assign m_14_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_15_io_y_3 = src1[32:30]; // @[MUL.scala 303:56]
  assign m_15_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_16_io_y_3 = src1[34:32]; // @[MUL.scala 303:56]
  assign m_16_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_17_io_y_3 = src1[36:34]; // @[MUL.scala 303:56]
  assign m_17_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_18_io_y_3 = src1[38:36]; // @[MUL.scala 303:56]
  assign m_18_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_19_io_y_3 = src1[40:38]; // @[MUL.scala 303:56]
  assign m_19_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_20_io_y_3 = src1[42:40]; // @[MUL.scala 303:56]
  assign m_20_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_21_io_y_3 = src1[44:42]; // @[MUL.scala 303:56]
  assign m_21_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_22_io_y_3 = src1[46:44]; // @[MUL.scala 303:56]
  assign m_22_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_23_io_y_3 = src1[48:46]; // @[MUL.scala 303:56]
  assign m_23_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_24_io_y_3 = src1[50:48]; // @[MUL.scala 303:56]
  assign m_24_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_25_io_y_3 = src1[52:50]; // @[MUL.scala 303:56]
  assign m_25_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_26_io_y_3 = src1[54:52]; // @[MUL.scala 303:56]
  assign m_26_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_27_io_y_3 = src1[56:54]; // @[MUL.scala 303:56]
  assign m_27_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_28_io_y_3 = src1[58:56]; // @[MUL.scala 303:56]
  assign m_28_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_29_io_y_3 = src1[60:58]; // @[MUL.scala 303:56]
  assign m_29_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_30_io_y_3 = src1[62:60]; // @[MUL.scala 303:56]
  assign m_30_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_31_io_y_3 = src1[64:62]; // @[MUL.scala 303:56]
  assign m_31_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_32_io_y_3 = src1[66:64]; // @[MUL.scala 303:56]
  assign m_32_io_x = {2'h0,io_in_bits_ctrl_data_src2}; // @[Cat.scala 31:58]
  assign m_33_io_in_0 = r; // @[MUL.scala 125:16]
  assign m_33_io_in_1 = r_1; // @[MUL.scala 126:16]
  assign m_34_io_in_0 = r_2; // @[MUL.scala 125:16]
  assign m_34_io_in_1 = r_3; // @[MUL.scala 126:16]
  assign m_35_io_x1 = r_4; // @[MUL.scala 103:13]
  assign m_35_io_x2 = r_5; // @[MUL.scala 104:13]
  assign m_35_io_x3 = r_6; // @[MUL.scala 105:13]
  assign m_36_io_x1 = r_7; // @[MUL.scala 103:13]
  assign m_36_io_x2 = r_8; // @[MUL.scala 104:13]
  assign m_36_io_x3 = r_9; // @[MUL.scala 105:13]
  assign m_37_io_x1 = r_10; // @[MUL.scala 103:13]
  assign m_37_io_x2 = r_11; // @[MUL.scala 104:13]
  assign m_37_io_x3 = r_12; // @[MUL.scala 105:13]
  assign m_38_io_x1 = r_14; // @[MUL.scala 103:13]
  assign m_38_io_x2 = r_15; // @[MUL.scala 104:13]
  assign m_38_io_x3 = r_16; // @[MUL.scala 105:13]
  assign m_39_io_x1 = r_18; // @[MUL.scala 103:13]
  assign m_39_io_x2 = r_19; // @[MUL.scala 104:13]
  assign m_39_io_x3 = r_20; // @[MUL.scala 105:13]
  assign m_40_io_in_0 = r_21; // @[MUL.scala 125:16]
  assign m_40_io_in_1 = r_22; // @[MUL.scala 126:16]
  assign m_41_io_x1 = r_23; // @[MUL.scala 103:13]
  assign m_41_io_x2 = r_24; // @[MUL.scala 104:13]
  assign m_41_io_x3 = r_25; // @[MUL.scala 105:13]
  assign m_42_io_in_0 = r_26; // @[MUL.scala 125:16]
  assign m_42_io_in_1 = r_27; // @[MUL.scala 126:16]
  assign m_43_io_x1 = r_28; // @[MUL.scala 103:13]
  assign m_43_io_x2 = r_29; // @[MUL.scala 104:13]
  assign m_43_io_x3 = r_30; // @[MUL.scala 105:13]
  assign m_44_io_x1 = r_31; // @[MUL.scala 103:13]
  assign m_44_io_x2 = r_32; // @[MUL.scala 104:13]
  assign m_44_io_x3 = r_33; // @[MUL.scala 105:13]
  assign m_45_io_x1 = r_34; // @[MUL.scala 103:13]
  assign m_45_io_x2 = r_35; // @[MUL.scala 104:13]
  assign m_45_io_x3 = r_36; // @[MUL.scala 105:13]
  assign m_46_io_x1 = r_37; // @[MUL.scala 103:13]
  assign m_46_io_x2 = r_38; // @[MUL.scala 104:13]
  assign m_46_io_x3 = r_39; // @[MUL.scala 105:13]
  assign m_47_io_x1 = r_40; // @[MUL.scala 103:13]
  assign m_47_io_x2 = r_41; // @[MUL.scala 104:13]
  assign m_47_io_x3 = r_42; // @[MUL.scala 105:13]
  assign m_48_io_x1 = r_43; // @[MUL.scala 103:13]
  assign m_48_io_x2 = r_44; // @[MUL.scala 104:13]
  assign m_48_io_x3 = r_45; // @[MUL.scala 105:13]
  assign m_49_io_x1 = r_47; // @[MUL.scala 103:13]
  assign m_49_io_x2 = r_48; // @[MUL.scala 104:13]
  assign m_49_io_x3 = r_49; // @[MUL.scala 105:13]
  assign m_50_io_x1 = r_50; // @[MUL.scala 103:13]
  assign m_50_io_x2 = r_51; // @[MUL.scala 104:13]
  assign m_50_io_x3 = r_52; // @[MUL.scala 105:13]
  assign m_51_io_x1 = r_54; // @[MUL.scala 103:13]
  assign m_51_io_x2 = r_55; // @[MUL.scala 104:13]
  assign m_51_io_x3 = r_56; // @[MUL.scala 105:13]
  assign m_52_io_x1 = r_57; // @[MUL.scala 103:13]
  assign m_52_io_x2 = r_58; // @[MUL.scala 104:13]
  assign m_52_io_x3 = r_59; // @[MUL.scala 105:13]
  assign m_53_io_in_0 = r_60; // @[MUL.scala 125:16]
  assign m_53_io_in_1 = r_61; // @[MUL.scala 126:16]
  assign m_54_io_x1 = r_62; // @[MUL.scala 103:13]
  assign m_54_io_x2 = r_63; // @[MUL.scala 104:13]
  assign m_54_io_x3 = r_64; // @[MUL.scala 105:13]
  assign m_55_io_x1 = r_65; // @[MUL.scala 103:13]
  assign m_55_io_x2 = r_66; // @[MUL.scala 104:13]
  assign m_55_io_x3 = r_67; // @[MUL.scala 105:13]
  assign m_56_io_in_0 = r_68; // @[MUL.scala 125:16]
  assign m_56_io_in_1 = r_69; // @[MUL.scala 126:16]
  assign m_57_io_x1 = r_70; // @[MUL.scala 103:13]
  assign m_57_io_x2 = r_71; // @[MUL.scala 104:13]
  assign m_57_io_x3 = r_72; // @[MUL.scala 105:13]
  assign m_58_io_x1 = r_73; // @[MUL.scala 103:13]
  assign m_58_io_x2 = r_74; // @[MUL.scala 104:13]
  assign m_58_io_x3 = r_75; // @[MUL.scala 105:13]
  assign m_59_io_x1 = r_76; // @[MUL.scala 103:13]
  assign m_59_io_x2 = r_77; // @[MUL.scala 104:13]
  assign m_59_io_x3 = r_78; // @[MUL.scala 105:13]
  assign m_60_io_x1 = r_79; // @[MUL.scala 103:13]
  assign m_60_io_x2 = r_80; // @[MUL.scala 104:13]
  assign m_60_io_x3 = r_81; // @[MUL.scala 105:13]
  assign m_61_io_x1 = r_82; // @[MUL.scala 103:13]
  assign m_61_io_x2 = r_83; // @[MUL.scala 104:13]
  assign m_61_io_x3 = r_84; // @[MUL.scala 105:13]
  assign m_62_io_x1 = r_85; // @[MUL.scala 103:13]
  assign m_62_io_x2 = r_86; // @[MUL.scala 104:13]
  assign m_62_io_x3 = r_87; // @[MUL.scala 105:13]
  assign m_63_io_x1 = r_88; // @[MUL.scala 103:13]
  assign m_63_io_x2 = r_89; // @[MUL.scala 104:13]
  assign m_63_io_x3 = r_90; // @[MUL.scala 105:13]
  assign m_64_io_x1 = r_91; // @[MUL.scala 103:13]
  assign m_64_io_x2 = r_92; // @[MUL.scala 104:13]
  assign m_64_io_x3 = r_93; // @[MUL.scala 105:13]
  assign m_65_io_x1 = r_94; // @[MUL.scala 103:13]
  assign m_65_io_x2 = r_95; // @[MUL.scala 104:13]
  assign m_65_io_x3 = r_96; // @[MUL.scala 105:13]
  assign m_66_io_x1 = r_98; // @[MUL.scala 103:13]
  assign m_66_io_x2 = r_99; // @[MUL.scala 104:13]
  assign m_66_io_x3 = r_100; // @[MUL.scala 105:13]
  assign m_67_io_x1 = r_101; // @[MUL.scala 103:13]
  assign m_67_io_x2 = r_102; // @[MUL.scala 104:13]
  assign m_67_io_x3 = r_103; // @[MUL.scala 105:13]
  assign m_68_io_x1 = r_104; // @[MUL.scala 103:13]
  assign m_68_io_x2 = r_105; // @[MUL.scala 104:13]
  assign m_68_io_x3 = r_106; // @[MUL.scala 105:13]
  assign m_69_io_x1 = r_108; // @[MUL.scala 103:13]
  assign m_69_io_x2 = r_109; // @[MUL.scala 104:13]
  assign m_69_io_x3 = r_110; // @[MUL.scala 105:13]
  assign m_70_io_x1 = r_111; // @[MUL.scala 103:13]
  assign m_70_io_x2 = r_112; // @[MUL.scala 104:13]
  assign m_70_io_x3 = r_113; // @[MUL.scala 105:13]
  assign m_71_io_x1 = r_114; // @[MUL.scala 103:13]
  assign m_71_io_x2 = r_115; // @[MUL.scala 104:13]
  assign m_71_io_x3 = r_116; // @[MUL.scala 105:13]
  assign m_72_io_in_0 = r_117; // @[MUL.scala 125:16]
  assign m_72_io_in_1 = r_118; // @[MUL.scala 126:16]
  assign m_73_io_x1 = r_119; // @[MUL.scala 103:13]
  assign m_73_io_x2 = r_120; // @[MUL.scala 104:13]
  assign m_73_io_x3 = r_121; // @[MUL.scala 105:13]
  assign m_74_io_x1 = r_122; // @[MUL.scala 103:13]
  assign m_74_io_x2 = r_123; // @[MUL.scala 104:13]
  assign m_74_io_x3 = r_124; // @[MUL.scala 105:13]
  assign m_75_io_x1 = r_125; // @[MUL.scala 103:13]
  assign m_75_io_x2 = r_126; // @[MUL.scala 104:13]
  assign m_75_io_x3 = r_127; // @[MUL.scala 105:13]
  assign m_76_io_in_0 = r_128; // @[MUL.scala 125:16]
  assign m_76_io_in_1 = r_129; // @[MUL.scala 126:16]
  assign m_77_io_x1 = r_130; // @[MUL.scala 103:13]
  assign m_77_io_x2 = r_131; // @[MUL.scala 104:13]
  assign m_77_io_x3 = r_132; // @[MUL.scala 105:13]
  assign m_78_io_x1 = r_133; // @[MUL.scala 103:13]
  assign m_78_io_x2 = r_134; // @[MUL.scala 104:13]
  assign m_78_io_x3 = r_135; // @[MUL.scala 105:13]
  assign m_79_io_x1 = r_136; // @[MUL.scala 103:13]
  assign m_79_io_x2 = r_137; // @[MUL.scala 104:13]
  assign m_79_io_x3 = r_138; // @[MUL.scala 105:13]
  assign m_80_io_x1 = r_139; // @[MUL.scala 103:13]
  assign m_80_io_x2 = r_140; // @[MUL.scala 104:13]
  assign m_80_io_x3 = r_141; // @[MUL.scala 105:13]
  assign m_81_io_x1 = r_142; // @[MUL.scala 103:13]
  assign m_81_io_x2 = r_143; // @[MUL.scala 104:13]
  assign m_81_io_x3 = r_144; // @[MUL.scala 105:13]
  assign m_82_io_x1 = r_145; // @[MUL.scala 103:13]
  assign m_82_io_x2 = r_146; // @[MUL.scala 104:13]
  assign m_82_io_x3 = r_147; // @[MUL.scala 105:13]
  assign m_83_io_x1 = r_148; // @[MUL.scala 103:13]
  assign m_83_io_x2 = r_149; // @[MUL.scala 104:13]
  assign m_83_io_x3 = r_150; // @[MUL.scala 105:13]
  assign m_84_io_x1 = r_151; // @[MUL.scala 103:13]
  assign m_84_io_x2 = r_152; // @[MUL.scala 104:13]
  assign m_84_io_x3 = r_153; // @[MUL.scala 105:13]
  assign m_85_io_x1 = r_154; // @[MUL.scala 103:13]
  assign m_85_io_x2 = r_155; // @[MUL.scala 104:13]
  assign m_85_io_x3 = r_156; // @[MUL.scala 105:13]
  assign m_86_io_x1 = r_157; // @[MUL.scala 103:13]
  assign m_86_io_x2 = r_158; // @[MUL.scala 104:13]
  assign m_86_io_x3 = r_159; // @[MUL.scala 105:13]
  assign m_87_io_x1 = r_160; // @[MUL.scala 103:13]
  assign m_87_io_x2 = r_161; // @[MUL.scala 104:13]
  assign m_87_io_x3 = r_162; // @[MUL.scala 105:13]
  assign m_88_io_x1 = r_163; // @[MUL.scala 103:13]
  assign m_88_io_x2 = r_164; // @[MUL.scala 104:13]
  assign m_88_io_x3 = r_165; // @[MUL.scala 105:13]
  assign m_89_io_x1 = r_167; // @[MUL.scala 103:13]
  assign m_89_io_x2 = r_168; // @[MUL.scala 104:13]
  assign m_89_io_x3 = r_169; // @[MUL.scala 105:13]
  assign m_90_io_x1 = r_170; // @[MUL.scala 103:13]
  assign m_90_io_x2 = r_171; // @[MUL.scala 104:13]
  assign m_90_io_x3 = r_172; // @[MUL.scala 105:13]
  assign m_91_io_x1 = r_173; // @[MUL.scala 103:13]
  assign m_91_io_x2 = r_174; // @[MUL.scala 104:13]
  assign m_91_io_x3 = r_175; // @[MUL.scala 105:13]
  assign m_92_io_x1 = r_176; // @[MUL.scala 103:13]
  assign m_92_io_x2 = r_177; // @[MUL.scala 104:13]
  assign m_92_io_x3 = r_178; // @[MUL.scala 105:13]
  assign m_93_io_x1 = r_180; // @[MUL.scala 103:13]
  assign m_93_io_x2 = r_181; // @[MUL.scala 104:13]
  assign m_93_io_x3 = r_182; // @[MUL.scala 105:13]
  assign m_94_io_x1 = r_183; // @[MUL.scala 103:13]
  assign m_94_io_x2 = r_184; // @[MUL.scala 104:13]
  assign m_94_io_x3 = r_185; // @[MUL.scala 105:13]
  assign m_95_io_x1 = r_186; // @[MUL.scala 103:13]
  assign m_95_io_x2 = r_187; // @[MUL.scala 104:13]
  assign m_95_io_x3 = r_188; // @[MUL.scala 105:13]
  assign m_96_io_x1 = r_189; // @[MUL.scala 103:13]
  assign m_96_io_x2 = r_190; // @[MUL.scala 104:13]
  assign m_96_io_x3 = r_191; // @[MUL.scala 105:13]
  assign m_97_io_in_0 = r_192; // @[MUL.scala 125:16]
  assign m_97_io_in_1 = r_193; // @[MUL.scala 126:16]
  assign m_98_io_x1 = r_194; // @[MUL.scala 103:13]
  assign m_98_io_x2 = r_195; // @[MUL.scala 104:13]
  assign m_98_io_x3 = r_196; // @[MUL.scala 105:13]
  assign m_99_io_x1 = r_197; // @[MUL.scala 103:13]
  assign m_99_io_x2 = r_198; // @[MUL.scala 104:13]
  assign m_99_io_x3 = r_199; // @[MUL.scala 105:13]
  assign m_100_io_x1 = r_200; // @[MUL.scala 103:13]
  assign m_100_io_x2 = r_201; // @[MUL.scala 104:13]
  assign m_100_io_x3 = r_202; // @[MUL.scala 105:13]
  assign m_101_io_x1 = r_203; // @[MUL.scala 103:13]
  assign m_101_io_x2 = r_204; // @[MUL.scala 104:13]
  assign m_101_io_x3 = r_205; // @[MUL.scala 105:13]
  assign m_102_io_in_0 = r_206; // @[MUL.scala 125:16]
  assign m_102_io_in_1 = r_207; // @[MUL.scala 126:16]
  assign m_103_io_x1 = r_208; // @[MUL.scala 103:13]
  assign m_103_io_x2 = r_209; // @[MUL.scala 104:13]
  assign m_103_io_x3 = r_210; // @[MUL.scala 105:13]
  assign m_104_io_x1 = r_211; // @[MUL.scala 103:13]
  assign m_104_io_x2 = r_212; // @[MUL.scala 104:13]
  assign m_104_io_x3 = r_213; // @[MUL.scala 105:13]
  assign m_105_io_x1 = r_214; // @[MUL.scala 103:13]
  assign m_105_io_x2 = r_215; // @[MUL.scala 104:13]
  assign m_105_io_x3 = r_216; // @[MUL.scala 105:13]
  assign m_106_io_x1 = r_217; // @[MUL.scala 103:13]
  assign m_106_io_x2 = r_218; // @[MUL.scala 104:13]
  assign m_106_io_x3 = r_219; // @[MUL.scala 105:13]
  assign m_107_io_x1 = r_220; // @[MUL.scala 103:13]
  assign m_107_io_x2 = r_221; // @[MUL.scala 104:13]
  assign m_107_io_x3 = r_222; // @[MUL.scala 105:13]
  assign m_108_io_x1 = r_223; // @[MUL.scala 103:13]
  assign m_108_io_x2 = r_224; // @[MUL.scala 104:13]
  assign m_108_io_x3 = r_225; // @[MUL.scala 105:13]
  assign m_109_io_x1 = r_226; // @[MUL.scala 103:13]
  assign m_109_io_x2 = r_227; // @[MUL.scala 104:13]
  assign m_109_io_x3 = r_228; // @[MUL.scala 105:13]
  assign m_110_io_x1 = r_229; // @[MUL.scala 103:13]
  assign m_110_io_x2 = r_230; // @[MUL.scala 104:13]
  assign m_110_io_x3 = r_231; // @[MUL.scala 105:13]
  assign m_111_io_x1 = r_232; // @[MUL.scala 103:13]
  assign m_111_io_x2 = r_233; // @[MUL.scala 104:13]
  assign m_111_io_x3 = r_234; // @[MUL.scala 105:13]
  assign m_112_io_x1 = r_235; // @[MUL.scala 103:13]
  assign m_112_io_x2 = r_236; // @[MUL.scala 104:13]
  assign m_112_io_x3 = r_237; // @[MUL.scala 105:13]
  assign m_113_io_x1 = r_238; // @[MUL.scala 103:13]
  assign m_113_io_x2 = r_239; // @[MUL.scala 104:13]
  assign m_113_io_x3 = r_240; // @[MUL.scala 105:13]
  assign m_114_io_x1 = r_241; // @[MUL.scala 103:13]
  assign m_114_io_x2 = r_242; // @[MUL.scala 104:13]
  assign m_114_io_x3 = r_243; // @[MUL.scala 105:13]
  assign m_115_io_x1 = r_244; // @[MUL.scala 103:13]
  assign m_115_io_x2 = r_245; // @[MUL.scala 104:13]
  assign m_115_io_x3 = r_246; // @[MUL.scala 105:13]
  assign m_116_io_x1 = r_247; // @[MUL.scala 103:13]
  assign m_116_io_x2 = r_248; // @[MUL.scala 104:13]
  assign m_116_io_x3 = r_249; // @[MUL.scala 105:13]
  assign m_117_io_x1 = r_250; // @[MUL.scala 103:13]
  assign m_117_io_x2 = r_251; // @[MUL.scala 104:13]
  assign m_117_io_x3 = r_252; // @[MUL.scala 105:13]
  assign m_118_io_x1 = r_254; // @[MUL.scala 103:13]
  assign m_118_io_x2 = r_255; // @[MUL.scala 104:13]
  assign m_118_io_x3 = r_256; // @[MUL.scala 105:13]
  assign m_119_io_x1 = r_257; // @[MUL.scala 103:13]
  assign m_119_io_x2 = r_258; // @[MUL.scala 104:13]
  assign m_119_io_x3 = r_259; // @[MUL.scala 105:13]
  assign m_120_io_x1 = r_260; // @[MUL.scala 103:13]
  assign m_120_io_x2 = r_261; // @[MUL.scala 104:13]
  assign m_120_io_x3 = r_262; // @[MUL.scala 105:13]
  assign m_121_io_x1 = r_263; // @[MUL.scala 103:13]
  assign m_121_io_x2 = r_264; // @[MUL.scala 104:13]
  assign m_121_io_x3 = r_265; // @[MUL.scala 105:13]
  assign m_122_io_x1 = r_266; // @[MUL.scala 103:13]
  assign m_122_io_x2 = r_267; // @[MUL.scala 104:13]
  assign m_122_io_x3 = r_268; // @[MUL.scala 105:13]
  assign m_123_io_x1 = r_270; // @[MUL.scala 103:13]
  assign m_123_io_x2 = r_271; // @[MUL.scala 104:13]
  assign m_123_io_x3 = r_272; // @[MUL.scala 105:13]
  assign m_124_io_x1 = r_273; // @[MUL.scala 103:13]
  assign m_124_io_x2 = r_274; // @[MUL.scala 104:13]
  assign m_124_io_x3 = r_275; // @[MUL.scala 105:13]
  assign m_125_io_x1 = r_276; // @[MUL.scala 103:13]
  assign m_125_io_x2 = r_277; // @[MUL.scala 104:13]
  assign m_125_io_x3 = r_278; // @[MUL.scala 105:13]
  assign m_126_io_x1 = r_279; // @[MUL.scala 103:13]
  assign m_126_io_x2 = r_280; // @[MUL.scala 104:13]
  assign m_126_io_x3 = r_281; // @[MUL.scala 105:13]
  assign m_127_io_x1 = r_282; // @[MUL.scala 103:13]
  assign m_127_io_x2 = r_283; // @[MUL.scala 104:13]
  assign m_127_io_x3 = r_284; // @[MUL.scala 105:13]
  assign m_128_io_in_0 = r_285; // @[MUL.scala 125:16]
  assign m_128_io_in_1 = r_286; // @[MUL.scala 126:16]
  assign m_129_io_x1 = r_287; // @[MUL.scala 103:13]
  assign m_129_io_x2 = r_288; // @[MUL.scala 104:13]
  assign m_129_io_x3 = r_289; // @[MUL.scala 105:13]
  assign m_130_io_x1 = r_290; // @[MUL.scala 103:13]
  assign m_130_io_x2 = r_291; // @[MUL.scala 104:13]
  assign m_130_io_x3 = r_292; // @[MUL.scala 105:13]
  assign m_131_io_x1 = r_293; // @[MUL.scala 103:13]
  assign m_131_io_x2 = r_294; // @[MUL.scala 104:13]
  assign m_131_io_x3 = r_295; // @[MUL.scala 105:13]
  assign m_132_io_x1 = r_296; // @[MUL.scala 103:13]
  assign m_132_io_x2 = r_297; // @[MUL.scala 104:13]
  assign m_132_io_x3 = r_298; // @[MUL.scala 105:13]
  assign m_133_io_x1 = r_299; // @[MUL.scala 103:13]
  assign m_133_io_x2 = r_300; // @[MUL.scala 104:13]
  assign m_133_io_x3 = r_301; // @[MUL.scala 105:13]
  assign m_134_io_in_0 = r_302; // @[MUL.scala 125:16]
  assign m_134_io_in_1 = r_303; // @[MUL.scala 126:16]
  assign m_135_io_x1 = r_304; // @[MUL.scala 103:13]
  assign m_135_io_x2 = r_305; // @[MUL.scala 104:13]
  assign m_135_io_x3 = r_306; // @[MUL.scala 105:13]
  assign m_136_io_x1 = r_307; // @[MUL.scala 103:13]
  assign m_136_io_x2 = r_308; // @[MUL.scala 104:13]
  assign m_136_io_x3 = r_309; // @[MUL.scala 105:13]
  assign m_137_io_x1 = r_310; // @[MUL.scala 103:13]
  assign m_137_io_x2 = r_311; // @[MUL.scala 104:13]
  assign m_137_io_x3 = r_312; // @[MUL.scala 105:13]
  assign m_138_io_x1 = r_313; // @[MUL.scala 103:13]
  assign m_138_io_x2 = r_314; // @[MUL.scala 104:13]
  assign m_138_io_x3 = r_315; // @[MUL.scala 105:13]
  assign m_139_io_x1 = r_316; // @[MUL.scala 103:13]
  assign m_139_io_x2 = r_317; // @[MUL.scala 104:13]
  assign m_139_io_x3 = r_318; // @[MUL.scala 105:13]
  assign m_140_io_x1 = r_319; // @[MUL.scala 103:13]
  assign m_140_io_x2 = r_320; // @[MUL.scala 104:13]
  assign m_140_io_x3 = r_321; // @[MUL.scala 105:13]
  assign m_141_io_x1 = r_322; // @[MUL.scala 103:13]
  assign m_141_io_x2 = r_323; // @[MUL.scala 104:13]
  assign m_141_io_x3 = r_324; // @[MUL.scala 105:13]
  assign m_142_io_x1 = r_325; // @[MUL.scala 103:13]
  assign m_142_io_x2 = r_326; // @[MUL.scala 104:13]
  assign m_142_io_x3 = r_327; // @[MUL.scala 105:13]
  assign m_143_io_x1 = r_328; // @[MUL.scala 103:13]
  assign m_143_io_x2 = r_329; // @[MUL.scala 104:13]
  assign m_143_io_x3 = r_330; // @[MUL.scala 105:13]
  assign m_144_io_x1 = r_331; // @[MUL.scala 103:13]
  assign m_144_io_x2 = r_332; // @[MUL.scala 104:13]
  assign m_144_io_x3 = r_333; // @[MUL.scala 105:13]
  assign m_145_io_x1 = r_334; // @[MUL.scala 103:13]
  assign m_145_io_x2 = r_335; // @[MUL.scala 104:13]
  assign m_145_io_x3 = r_336; // @[MUL.scala 105:13]
  assign m_146_io_x1 = r_337; // @[MUL.scala 103:13]
  assign m_146_io_x2 = r_338; // @[MUL.scala 104:13]
  assign m_146_io_x3 = r_339; // @[MUL.scala 105:13]
  assign m_147_io_x1 = r_340; // @[MUL.scala 103:13]
  assign m_147_io_x2 = r_341; // @[MUL.scala 104:13]
  assign m_147_io_x3 = r_342; // @[MUL.scala 105:13]
  assign m_148_io_x1 = r_343; // @[MUL.scala 103:13]
  assign m_148_io_x2 = r_344; // @[MUL.scala 104:13]
  assign m_148_io_x3 = r_345; // @[MUL.scala 105:13]
  assign m_149_io_x1 = r_346; // @[MUL.scala 103:13]
  assign m_149_io_x2 = r_347; // @[MUL.scala 104:13]
  assign m_149_io_x3 = r_348; // @[MUL.scala 105:13]
  assign m_150_io_x1 = r_349; // @[MUL.scala 103:13]
  assign m_150_io_x2 = r_350; // @[MUL.scala 104:13]
  assign m_150_io_x3 = r_351; // @[MUL.scala 105:13]
  assign m_151_io_x1 = r_352; // @[MUL.scala 103:13]
  assign m_151_io_x2 = r_353; // @[MUL.scala 104:13]
  assign m_151_io_x3 = r_354; // @[MUL.scala 105:13]
  assign m_152_io_x1 = r_355; // @[MUL.scala 103:13]
  assign m_152_io_x2 = r_356; // @[MUL.scala 104:13]
  assign m_152_io_x3 = r_357; // @[MUL.scala 105:13]
  assign m_153_io_x1 = r_359; // @[MUL.scala 103:13]
  assign m_153_io_x2 = r_360; // @[MUL.scala 104:13]
  assign m_153_io_x3 = r_361; // @[MUL.scala 105:13]
  assign m_154_io_x1 = r_362; // @[MUL.scala 103:13]
  assign m_154_io_x2 = r_363; // @[MUL.scala 104:13]
  assign m_154_io_x3 = r_364; // @[MUL.scala 105:13]
  assign m_155_io_x1 = r_365; // @[MUL.scala 103:13]
  assign m_155_io_x2 = r_366; // @[MUL.scala 104:13]
  assign m_155_io_x3 = r_367; // @[MUL.scala 105:13]
  assign m_156_io_x1 = r_368; // @[MUL.scala 103:13]
  assign m_156_io_x2 = r_369; // @[MUL.scala 104:13]
  assign m_156_io_x3 = r_370; // @[MUL.scala 105:13]
  assign m_157_io_x1 = r_371; // @[MUL.scala 103:13]
  assign m_157_io_x2 = r_372; // @[MUL.scala 104:13]
  assign m_157_io_x3 = r_373; // @[MUL.scala 105:13]
  assign m_158_io_x1 = r_374; // @[MUL.scala 103:13]
  assign m_158_io_x2 = r_375; // @[MUL.scala 104:13]
  assign m_158_io_x3 = r_376; // @[MUL.scala 105:13]
  assign m_159_io_x1 = r_378; // @[MUL.scala 103:13]
  assign m_159_io_x2 = r_379; // @[MUL.scala 104:13]
  assign m_159_io_x3 = r_380; // @[MUL.scala 105:13]
  assign m_160_io_x1 = r_381; // @[MUL.scala 103:13]
  assign m_160_io_x2 = r_382; // @[MUL.scala 104:13]
  assign m_160_io_x3 = r_383; // @[MUL.scala 105:13]
  assign m_161_io_x1 = r_384; // @[MUL.scala 103:13]
  assign m_161_io_x2 = r_385; // @[MUL.scala 104:13]
  assign m_161_io_x3 = r_386; // @[MUL.scala 105:13]
  assign m_162_io_x1 = r_387; // @[MUL.scala 103:13]
  assign m_162_io_x2 = r_388; // @[MUL.scala 104:13]
  assign m_162_io_x3 = r_389; // @[MUL.scala 105:13]
  assign m_163_io_x1 = r_390; // @[MUL.scala 103:13]
  assign m_163_io_x2 = r_391; // @[MUL.scala 104:13]
  assign m_163_io_x3 = r_392; // @[MUL.scala 105:13]
  assign m_164_io_x1 = r_393; // @[MUL.scala 103:13]
  assign m_164_io_x2 = r_394; // @[MUL.scala 104:13]
  assign m_164_io_x3 = r_395; // @[MUL.scala 105:13]
  assign m_165_io_in_0 = r_396; // @[MUL.scala 125:16]
  assign m_165_io_in_1 = r_397; // @[MUL.scala 126:16]
  assign m_166_io_x1 = r_398; // @[MUL.scala 103:13]
  assign m_166_io_x2 = r_399; // @[MUL.scala 104:13]
  assign m_166_io_x3 = r_400; // @[MUL.scala 105:13]
  assign m_167_io_x1 = r_401; // @[MUL.scala 103:13]
  assign m_167_io_x2 = r_402; // @[MUL.scala 104:13]
  assign m_167_io_x3 = r_403; // @[MUL.scala 105:13]
  assign m_168_io_x1 = r_404; // @[MUL.scala 103:13]
  assign m_168_io_x2 = r_405; // @[MUL.scala 104:13]
  assign m_168_io_x3 = r_406; // @[MUL.scala 105:13]
  assign m_169_io_x1 = r_407; // @[MUL.scala 103:13]
  assign m_169_io_x2 = r_408; // @[MUL.scala 104:13]
  assign m_169_io_x3 = r_409; // @[MUL.scala 105:13]
  assign m_170_io_x1 = r_410; // @[MUL.scala 103:13]
  assign m_170_io_x2 = r_411; // @[MUL.scala 104:13]
  assign m_170_io_x3 = r_412; // @[MUL.scala 105:13]
  assign m_171_io_x1 = r_413; // @[MUL.scala 103:13]
  assign m_171_io_x2 = r_414; // @[MUL.scala 104:13]
  assign m_171_io_x3 = r_415; // @[MUL.scala 105:13]
  assign m_172_io_in_0 = r_416; // @[MUL.scala 125:16]
  assign m_172_io_in_1 = r_417; // @[MUL.scala 126:16]
  assign m_173_io_x1 = r_418; // @[MUL.scala 103:13]
  assign m_173_io_x2 = r_419; // @[MUL.scala 104:13]
  assign m_173_io_x3 = r_420; // @[MUL.scala 105:13]
  assign m_174_io_x1 = r_421; // @[MUL.scala 103:13]
  assign m_174_io_x2 = r_422; // @[MUL.scala 104:13]
  assign m_174_io_x3 = r_423; // @[MUL.scala 105:13]
  assign m_175_io_x1 = r_424; // @[MUL.scala 103:13]
  assign m_175_io_x2 = r_425; // @[MUL.scala 104:13]
  assign m_175_io_x3 = r_426; // @[MUL.scala 105:13]
  assign m_176_io_x1 = r_427; // @[MUL.scala 103:13]
  assign m_176_io_x2 = r_428; // @[MUL.scala 104:13]
  assign m_176_io_x3 = r_429; // @[MUL.scala 105:13]
  assign m_177_io_x1 = r_430; // @[MUL.scala 103:13]
  assign m_177_io_x2 = r_431; // @[MUL.scala 104:13]
  assign m_177_io_x3 = r_432; // @[MUL.scala 105:13]
  assign m_178_io_x1 = r_433; // @[MUL.scala 103:13]
  assign m_178_io_x2 = r_434; // @[MUL.scala 104:13]
  assign m_178_io_x3 = r_435; // @[MUL.scala 105:13]
  assign m_179_io_x1 = r_436; // @[MUL.scala 103:13]
  assign m_179_io_x2 = r_437; // @[MUL.scala 104:13]
  assign m_179_io_x3 = r_438; // @[MUL.scala 105:13]
  assign m_180_io_x1 = r_439; // @[MUL.scala 103:13]
  assign m_180_io_x2 = r_440; // @[MUL.scala 104:13]
  assign m_180_io_x3 = r_441; // @[MUL.scala 105:13]
  assign m_181_io_x1 = r_442; // @[MUL.scala 103:13]
  assign m_181_io_x2 = r_443; // @[MUL.scala 104:13]
  assign m_181_io_x3 = r_444; // @[MUL.scala 105:13]
  assign m_182_io_x1 = r_445; // @[MUL.scala 103:13]
  assign m_182_io_x2 = r_446; // @[MUL.scala 104:13]
  assign m_182_io_x3 = r_447; // @[MUL.scala 105:13]
  assign m_183_io_x1 = r_448; // @[MUL.scala 103:13]
  assign m_183_io_x2 = r_449; // @[MUL.scala 104:13]
  assign m_183_io_x3 = r_450; // @[MUL.scala 105:13]
  assign m_184_io_x1 = r_451; // @[MUL.scala 103:13]
  assign m_184_io_x2 = r_452; // @[MUL.scala 104:13]
  assign m_184_io_x3 = r_453; // @[MUL.scala 105:13]
  assign m_185_io_x1 = r_454; // @[MUL.scala 103:13]
  assign m_185_io_x2 = r_455; // @[MUL.scala 104:13]
  assign m_185_io_x3 = r_456; // @[MUL.scala 105:13]
  assign m_186_io_x1 = r_457; // @[MUL.scala 103:13]
  assign m_186_io_x2 = r_458; // @[MUL.scala 104:13]
  assign m_186_io_x3 = r_459; // @[MUL.scala 105:13]
  assign m_187_io_x1 = r_460; // @[MUL.scala 103:13]
  assign m_187_io_x2 = r_461; // @[MUL.scala 104:13]
  assign m_187_io_x3 = r_462; // @[MUL.scala 105:13]
  assign m_188_io_x1 = r_463; // @[MUL.scala 103:13]
  assign m_188_io_x2 = r_464; // @[MUL.scala 104:13]
  assign m_188_io_x3 = r_465; // @[MUL.scala 105:13]
  assign m_189_io_x1 = r_466; // @[MUL.scala 103:13]
  assign m_189_io_x2 = r_467; // @[MUL.scala 104:13]
  assign m_189_io_x3 = r_468; // @[MUL.scala 105:13]
  assign m_190_io_x1 = r_469; // @[MUL.scala 103:13]
  assign m_190_io_x2 = r_470; // @[MUL.scala 104:13]
  assign m_190_io_x3 = r_471; // @[MUL.scala 105:13]
  assign m_191_io_x1 = r_472; // @[MUL.scala 103:13]
  assign m_191_io_x2 = r_473; // @[MUL.scala 104:13]
  assign m_191_io_x3 = r_474; // @[MUL.scala 105:13]
  assign m_192_io_x1 = r_475; // @[MUL.scala 103:13]
  assign m_192_io_x2 = r_476; // @[MUL.scala 104:13]
  assign m_192_io_x3 = r_477; // @[MUL.scala 105:13]
  assign m_193_io_x1 = r_478; // @[MUL.scala 103:13]
  assign m_193_io_x2 = r_479; // @[MUL.scala 104:13]
  assign m_193_io_x3 = r_480; // @[MUL.scala 105:13]
  assign m_194_io_x1 = r_482; // @[MUL.scala 103:13]
  assign m_194_io_x2 = r_483; // @[MUL.scala 104:13]
  assign m_194_io_x3 = r_484; // @[MUL.scala 105:13]
  assign m_195_io_x1 = r_485; // @[MUL.scala 103:13]
  assign m_195_io_x2 = r_486; // @[MUL.scala 104:13]
  assign m_195_io_x3 = r_487; // @[MUL.scala 105:13]
  assign m_196_io_x1 = r_488; // @[MUL.scala 103:13]
  assign m_196_io_x2 = r_489; // @[MUL.scala 104:13]
  assign m_196_io_x3 = r_490; // @[MUL.scala 105:13]
  assign m_197_io_x1 = r_491; // @[MUL.scala 103:13]
  assign m_197_io_x2 = r_492; // @[MUL.scala 104:13]
  assign m_197_io_x3 = r_493; // @[MUL.scala 105:13]
  assign m_198_io_x1 = r_494; // @[MUL.scala 103:13]
  assign m_198_io_x2 = r_495; // @[MUL.scala 104:13]
  assign m_198_io_x3 = r_496; // @[MUL.scala 105:13]
  assign m_199_io_x1 = r_497; // @[MUL.scala 103:13]
  assign m_199_io_x2 = r_498; // @[MUL.scala 104:13]
  assign m_199_io_x3 = r_499; // @[MUL.scala 105:13]
  assign m_200_io_x1 = r_500; // @[MUL.scala 103:13]
  assign m_200_io_x2 = r_501; // @[MUL.scala 104:13]
  assign m_200_io_x3 = r_502; // @[MUL.scala 105:13]
  assign m_201_io_x1 = r_504; // @[MUL.scala 103:13]
  assign m_201_io_x2 = r_505; // @[MUL.scala 104:13]
  assign m_201_io_x3 = r_506; // @[MUL.scala 105:13]
  assign m_202_io_x1 = r_507; // @[MUL.scala 103:13]
  assign m_202_io_x2 = r_508; // @[MUL.scala 104:13]
  assign m_202_io_x3 = r_509; // @[MUL.scala 105:13]
  assign m_203_io_x1 = r_510; // @[MUL.scala 103:13]
  assign m_203_io_x2 = r_511; // @[MUL.scala 104:13]
  assign m_203_io_x3 = r_512; // @[MUL.scala 105:13]
  assign m_204_io_x1 = r_513; // @[MUL.scala 103:13]
  assign m_204_io_x2 = r_514; // @[MUL.scala 104:13]
  assign m_204_io_x3 = r_515; // @[MUL.scala 105:13]
  assign m_205_io_x1 = r_516; // @[MUL.scala 103:13]
  assign m_205_io_x2 = r_517; // @[MUL.scala 104:13]
  assign m_205_io_x3 = r_518; // @[MUL.scala 105:13]
  assign m_206_io_x1 = r_519; // @[MUL.scala 103:13]
  assign m_206_io_x2 = r_520; // @[MUL.scala 104:13]
  assign m_206_io_x3 = r_521; // @[MUL.scala 105:13]
  assign m_207_io_x1 = r_522; // @[MUL.scala 103:13]
  assign m_207_io_x2 = r_523; // @[MUL.scala 104:13]
  assign m_207_io_x3 = r_524; // @[MUL.scala 105:13]
  assign m_208_io_in_0 = r_525; // @[MUL.scala 125:16]
  assign m_208_io_in_1 = r_526; // @[MUL.scala 126:16]
  assign m_209_io_x1 = r_527; // @[MUL.scala 103:13]
  assign m_209_io_x2 = r_528; // @[MUL.scala 104:13]
  assign m_209_io_x3 = r_529; // @[MUL.scala 105:13]
  assign m_210_io_x1 = r_530; // @[MUL.scala 103:13]
  assign m_210_io_x2 = r_531; // @[MUL.scala 104:13]
  assign m_210_io_x3 = r_532; // @[MUL.scala 105:13]
  assign m_211_io_x1 = r_533; // @[MUL.scala 103:13]
  assign m_211_io_x2 = r_534; // @[MUL.scala 104:13]
  assign m_211_io_x3 = r_535; // @[MUL.scala 105:13]
  assign m_212_io_x1 = r_536; // @[MUL.scala 103:13]
  assign m_212_io_x2 = r_537; // @[MUL.scala 104:13]
  assign m_212_io_x3 = r_538; // @[MUL.scala 105:13]
  assign m_213_io_x1 = r_539; // @[MUL.scala 103:13]
  assign m_213_io_x2 = r_540; // @[MUL.scala 104:13]
  assign m_213_io_x3 = r_541; // @[MUL.scala 105:13]
  assign m_214_io_x1 = r_542; // @[MUL.scala 103:13]
  assign m_214_io_x2 = r_543; // @[MUL.scala 104:13]
  assign m_214_io_x3 = r_544; // @[MUL.scala 105:13]
  assign m_215_io_x1 = r_545; // @[MUL.scala 103:13]
  assign m_215_io_x2 = r_546; // @[MUL.scala 104:13]
  assign m_215_io_x3 = r_547; // @[MUL.scala 105:13]
  assign m_216_io_in_0 = r_548; // @[MUL.scala 125:16]
  assign m_216_io_in_1 = r_549; // @[MUL.scala 126:16]
  assign m_217_io_x1 = r_550; // @[MUL.scala 103:13]
  assign m_217_io_x2 = r_551; // @[MUL.scala 104:13]
  assign m_217_io_x3 = r_552; // @[MUL.scala 105:13]
  assign m_218_io_x1 = r_553; // @[MUL.scala 103:13]
  assign m_218_io_x2 = r_554; // @[MUL.scala 104:13]
  assign m_218_io_x3 = r_555; // @[MUL.scala 105:13]
  assign m_219_io_x1 = r_556; // @[MUL.scala 103:13]
  assign m_219_io_x2 = r_557; // @[MUL.scala 104:13]
  assign m_219_io_x3 = r_558; // @[MUL.scala 105:13]
  assign m_220_io_x1 = r_559; // @[MUL.scala 103:13]
  assign m_220_io_x2 = r_560; // @[MUL.scala 104:13]
  assign m_220_io_x3 = r_561; // @[MUL.scala 105:13]
  assign m_221_io_x1 = r_562; // @[MUL.scala 103:13]
  assign m_221_io_x2 = r_563; // @[MUL.scala 104:13]
  assign m_221_io_x3 = r_564; // @[MUL.scala 105:13]
  assign m_222_io_x1 = r_565; // @[MUL.scala 103:13]
  assign m_222_io_x2 = r_566; // @[MUL.scala 104:13]
  assign m_222_io_x3 = r_567; // @[MUL.scala 105:13]
  assign m_223_io_x1 = r_568; // @[MUL.scala 103:13]
  assign m_223_io_x2 = r_569; // @[MUL.scala 104:13]
  assign m_223_io_x3 = r_570; // @[MUL.scala 105:13]
  assign m_224_io_x1 = r_571; // @[MUL.scala 103:13]
  assign m_224_io_x2 = r_572; // @[MUL.scala 104:13]
  assign m_224_io_x3 = r_573; // @[MUL.scala 105:13]
  assign m_225_io_x1 = r_574; // @[MUL.scala 103:13]
  assign m_225_io_x2 = r_575; // @[MUL.scala 104:13]
  assign m_225_io_x3 = r_576; // @[MUL.scala 105:13]
  assign m_226_io_x1 = r_577; // @[MUL.scala 103:13]
  assign m_226_io_x2 = r_578; // @[MUL.scala 104:13]
  assign m_226_io_x3 = r_579; // @[MUL.scala 105:13]
  assign m_227_io_x1 = r_580; // @[MUL.scala 103:13]
  assign m_227_io_x2 = r_581; // @[MUL.scala 104:13]
  assign m_227_io_x3 = r_582; // @[MUL.scala 105:13]
  assign m_228_io_x1 = r_583; // @[MUL.scala 103:13]
  assign m_228_io_x2 = r_584; // @[MUL.scala 104:13]
  assign m_228_io_x3 = r_585; // @[MUL.scala 105:13]
  assign m_229_io_x1 = r_586; // @[MUL.scala 103:13]
  assign m_229_io_x2 = r_587; // @[MUL.scala 104:13]
  assign m_229_io_x3 = r_588; // @[MUL.scala 105:13]
  assign m_230_io_x1 = r_589; // @[MUL.scala 103:13]
  assign m_230_io_x2 = r_590; // @[MUL.scala 104:13]
  assign m_230_io_x3 = r_591; // @[MUL.scala 105:13]
  assign m_231_io_x1 = r_592; // @[MUL.scala 103:13]
  assign m_231_io_x2 = r_593; // @[MUL.scala 104:13]
  assign m_231_io_x3 = r_594; // @[MUL.scala 105:13]
  assign m_232_io_x1 = r_595; // @[MUL.scala 103:13]
  assign m_232_io_x2 = r_596; // @[MUL.scala 104:13]
  assign m_232_io_x3 = r_597; // @[MUL.scala 105:13]
  assign m_233_io_x1 = r_598; // @[MUL.scala 103:13]
  assign m_233_io_x2 = r_599; // @[MUL.scala 104:13]
  assign m_233_io_x3 = r_600; // @[MUL.scala 105:13]
  assign m_234_io_x1 = r_601; // @[MUL.scala 103:13]
  assign m_234_io_x2 = r_602; // @[MUL.scala 104:13]
  assign m_234_io_x3 = r_603; // @[MUL.scala 105:13]
  assign m_235_io_x1 = r_604; // @[MUL.scala 103:13]
  assign m_235_io_x2 = r_605; // @[MUL.scala 104:13]
  assign m_235_io_x3 = r_606; // @[MUL.scala 105:13]
  assign m_236_io_x1 = r_607; // @[MUL.scala 103:13]
  assign m_236_io_x2 = r_608; // @[MUL.scala 104:13]
  assign m_236_io_x3 = r_609; // @[MUL.scala 105:13]
  assign m_237_io_x1 = r_610; // @[MUL.scala 103:13]
  assign m_237_io_x2 = r_611; // @[MUL.scala 104:13]
  assign m_237_io_x3 = r_612; // @[MUL.scala 105:13]
  assign m_238_io_x1 = r_613; // @[MUL.scala 103:13]
  assign m_238_io_x2 = r_614; // @[MUL.scala 104:13]
  assign m_238_io_x3 = r_615; // @[MUL.scala 105:13]
  assign m_239_io_x1 = r_616; // @[MUL.scala 103:13]
  assign m_239_io_x2 = r_617; // @[MUL.scala 104:13]
  assign m_239_io_x3 = r_618; // @[MUL.scala 105:13]
  assign m_240_io_x1 = r_619; // @[MUL.scala 103:13]
  assign m_240_io_x2 = r_620; // @[MUL.scala 104:13]
  assign m_240_io_x3 = r_621; // @[MUL.scala 105:13]
  assign m_241_io_x1 = r_623; // @[MUL.scala 103:13]
  assign m_241_io_x2 = r_624; // @[MUL.scala 104:13]
  assign m_241_io_x3 = r_625; // @[MUL.scala 105:13]
  assign m_242_io_x1 = r_626; // @[MUL.scala 103:13]
  assign m_242_io_x2 = r_627; // @[MUL.scala 104:13]
  assign m_242_io_x3 = r_628; // @[MUL.scala 105:13]
  assign m_243_io_x1 = r_629; // @[MUL.scala 103:13]
  assign m_243_io_x2 = r_630; // @[MUL.scala 104:13]
  assign m_243_io_x3 = r_631; // @[MUL.scala 105:13]
  assign m_244_io_x1 = r_632; // @[MUL.scala 103:13]
  assign m_244_io_x2 = r_633; // @[MUL.scala 104:13]
  assign m_244_io_x3 = r_634; // @[MUL.scala 105:13]
  assign m_245_io_x1 = r_635; // @[MUL.scala 103:13]
  assign m_245_io_x2 = r_636; // @[MUL.scala 104:13]
  assign m_245_io_x3 = r_637; // @[MUL.scala 105:13]
  assign m_246_io_x1 = r_638; // @[MUL.scala 103:13]
  assign m_246_io_x2 = r_639; // @[MUL.scala 104:13]
  assign m_246_io_x3 = r_640; // @[MUL.scala 105:13]
  assign m_247_io_x1 = r_641; // @[MUL.scala 103:13]
  assign m_247_io_x2 = r_642; // @[MUL.scala 104:13]
  assign m_247_io_x3 = r_643; // @[MUL.scala 105:13]
  assign m_248_io_x1 = r_644; // @[MUL.scala 103:13]
  assign m_248_io_x2 = r_645; // @[MUL.scala 104:13]
  assign m_248_io_x3 = r_646; // @[MUL.scala 105:13]
  assign m_249_io_x1 = r_648; // @[MUL.scala 103:13]
  assign m_249_io_x2 = r_649; // @[MUL.scala 104:13]
  assign m_249_io_x3 = r_650; // @[MUL.scala 105:13]
  assign m_250_io_x1 = r_651; // @[MUL.scala 103:13]
  assign m_250_io_x2 = r_652; // @[MUL.scala 104:13]
  assign m_250_io_x3 = r_653; // @[MUL.scala 105:13]
  assign m_251_io_x1 = r_654; // @[MUL.scala 103:13]
  assign m_251_io_x2 = r_655; // @[MUL.scala 104:13]
  assign m_251_io_x3 = r_656; // @[MUL.scala 105:13]
  assign m_252_io_x1 = r_657; // @[MUL.scala 103:13]
  assign m_252_io_x2 = r_658; // @[MUL.scala 104:13]
  assign m_252_io_x3 = r_659; // @[MUL.scala 105:13]
  assign m_253_io_x1 = r_660; // @[MUL.scala 103:13]
  assign m_253_io_x2 = r_661; // @[MUL.scala 104:13]
  assign m_253_io_x3 = r_662; // @[MUL.scala 105:13]
  assign m_254_io_x1 = r_663; // @[MUL.scala 103:13]
  assign m_254_io_x2 = r_664; // @[MUL.scala 104:13]
  assign m_254_io_x3 = r_665; // @[MUL.scala 105:13]
  assign m_255_io_x1 = r_666; // @[MUL.scala 103:13]
  assign m_255_io_x2 = r_667; // @[MUL.scala 104:13]
  assign m_255_io_x3 = r_668; // @[MUL.scala 105:13]
  assign m_256_io_x1 = r_669; // @[MUL.scala 103:13]
  assign m_256_io_x2 = r_670; // @[MUL.scala 104:13]
  assign m_256_io_x3 = r_671; // @[MUL.scala 105:13]
  assign m_257_io_in_0 = r_672; // @[MUL.scala 125:16]
  assign m_257_io_in_1 = r_673; // @[MUL.scala 126:16]
  assign m_258_io_x1 = r_674; // @[MUL.scala 103:13]
  assign m_258_io_x2 = r_675; // @[MUL.scala 104:13]
  assign m_258_io_x3 = r_676; // @[MUL.scala 105:13]
  assign m_259_io_x1 = r_677; // @[MUL.scala 103:13]
  assign m_259_io_x2 = r_678; // @[MUL.scala 104:13]
  assign m_259_io_x3 = r_679; // @[MUL.scala 105:13]
  assign m_260_io_x1 = r_680; // @[MUL.scala 103:13]
  assign m_260_io_x2 = r_681; // @[MUL.scala 104:13]
  assign m_260_io_x3 = r_682; // @[MUL.scala 105:13]
  assign m_261_io_x1 = r_683; // @[MUL.scala 103:13]
  assign m_261_io_x2 = r_684; // @[MUL.scala 104:13]
  assign m_261_io_x3 = r_685; // @[MUL.scala 105:13]
  assign m_262_io_x1 = r_686; // @[MUL.scala 103:13]
  assign m_262_io_x2 = r_687; // @[MUL.scala 104:13]
  assign m_262_io_x3 = r_688; // @[MUL.scala 105:13]
  assign m_263_io_x1 = r_689; // @[MUL.scala 103:13]
  assign m_263_io_x2 = r_690; // @[MUL.scala 104:13]
  assign m_263_io_x3 = r_691; // @[MUL.scala 105:13]
  assign m_264_io_x1 = r_692; // @[MUL.scala 103:13]
  assign m_264_io_x2 = r_693; // @[MUL.scala 104:13]
  assign m_264_io_x3 = r_694; // @[MUL.scala 105:13]
  assign m_265_io_x1 = r_695; // @[MUL.scala 103:13]
  assign m_265_io_x2 = r_696; // @[MUL.scala 104:13]
  assign m_265_io_x3 = r_697; // @[MUL.scala 105:13]
  assign m_266_io_in_0 = r_698; // @[MUL.scala 125:16]
  assign m_266_io_in_1 = r_699; // @[MUL.scala 126:16]
  assign m_267_io_x1 = r_700; // @[MUL.scala 103:13]
  assign m_267_io_x2 = r_701; // @[MUL.scala 104:13]
  assign m_267_io_x3 = r_702; // @[MUL.scala 105:13]
  assign m_268_io_x1 = r_703; // @[MUL.scala 103:13]
  assign m_268_io_x2 = r_704; // @[MUL.scala 104:13]
  assign m_268_io_x3 = r_705; // @[MUL.scala 105:13]
  assign m_269_io_x1 = r_706; // @[MUL.scala 103:13]
  assign m_269_io_x2 = r_707; // @[MUL.scala 104:13]
  assign m_269_io_x3 = r_708; // @[MUL.scala 105:13]
  assign m_270_io_x1 = r_709; // @[MUL.scala 103:13]
  assign m_270_io_x2 = r_710; // @[MUL.scala 104:13]
  assign m_270_io_x3 = r_711; // @[MUL.scala 105:13]
  assign m_271_io_x1 = r_712; // @[MUL.scala 103:13]
  assign m_271_io_x2 = r_713; // @[MUL.scala 104:13]
  assign m_271_io_x3 = r_714; // @[MUL.scala 105:13]
  assign m_272_io_x1 = r_715; // @[MUL.scala 103:13]
  assign m_272_io_x2 = r_716; // @[MUL.scala 104:13]
  assign m_272_io_x3 = r_717; // @[MUL.scala 105:13]
  assign m_273_io_x1 = r_718; // @[MUL.scala 103:13]
  assign m_273_io_x2 = r_719; // @[MUL.scala 104:13]
  assign m_273_io_x3 = r_720; // @[MUL.scala 105:13]
  assign m_274_io_x1 = r_721; // @[MUL.scala 103:13]
  assign m_274_io_x2 = r_722; // @[MUL.scala 104:13]
  assign m_274_io_x3 = r_723; // @[MUL.scala 105:13]
  assign m_275_io_x1 = r_724; // @[MUL.scala 103:13]
  assign m_275_io_x2 = r_725; // @[MUL.scala 104:13]
  assign m_275_io_x3 = r_726; // @[MUL.scala 105:13]
  assign m_276_io_x1 = r_727; // @[MUL.scala 103:13]
  assign m_276_io_x2 = r_728; // @[MUL.scala 104:13]
  assign m_276_io_x3 = r_729; // @[MUL.scala 105:13]
  assign m_277_io_x1 = r_730; // @[MUL.scala 103:13]
  assign m_277_io_x2 = r_731; // @[MUL.scala 104:13]
  assign m_277_io_x3 = r_732; // @[MUL.scala 105:13]
  assign m_278_io_x1 = r_733; // @[MUL.scala 103:13]
  assign m_278_io_x2 = r_734; // @[MUL.scala 104:13]
  assign m_278_io_x3 = r_735; // @[MUL.scala 105:13]
  assign m_279_io_x1 = r_736; // @[MUL.scala 103:13]
  assign m_279_io_x2 = r_737; // @[MUL.scala 104:13]
  assign m_279_io_x3 = r_738; // @[MUL.scala 105:13]
  assign m_280_io_x1 = r_739; // @[MUL.scala 103:13]
  assign m_280_io_x2 = r_740; // @[MUL.scala 104:13]
  assign m_280_io_x3 = r_741; // @[MUL.scala 105:13]
  assign m_281_io_x1 = r_742; // @[MUL.scala 103:13]
  assign m_281_io_x2 = r_743; // @[MUL.scala 104:13]
  assign m_281_io_x3 = r_744; // @[MUL.scala 105:13]
  assign m_282_io_x1 = r_745; // @[MUL.scala 103:13]
  assign m_282_io_x2 = r_746; // @[MUL.scala 104:13]
  assign m_282_io_x3 = r_747; // @[MUL.scala 105:13]
  assign m_283_io_x1 = r_748; // @[MUL.scala 103:13]
  assign m_283_io_x2 = r_749; // @[MUL.scala 104:13]
  assign m_283_io_x3 = r_750; // @[MUL.scala 105:13]
  assign m_284_io_x1 = r_751; // @[MUL.scala 103:13]
  assign m_284_io_x2 = r_752; // @[MUL.scala 104:13]
  assign m_284_io_x3 = r_753; // @[MUL.scala 105:13]
  assign m_285_io_x1 = r_754; // @[MUL.scala 103:13]
  assign m_285_io_x2 = r_755; // @[MUL.scala 104:13]
  assign m_285_io_x3 = r_756; // @[MUL.scala 105:13]
  assign m_286_io_x1 = r_757; // @[MUL.scala 103:13]
  assign m_286_io_x2 = r_758; // @[MUL.scala 104:13]
  assign m_286_io_x3 = r_759; // @[MUL.scala 105:13]
  assign m_287_io_x1 = r_760; // @[MUL.scala 103:13]
  assign m_287_io_x2 = r_761; // @[MUL.scala 104:13]
  assign m_287_io_x3 = r_762; // @[MUL.scala 105:13]
  assign m_288_io_x1 = r_763; // @[MUL.scala 103:13]
  assign m_288_io_x2 = r_764; // @[MUL.scala 104:13]
  assign m_288_io_x3 = r_765; // @[MUL.scala 105:13]
  assign m_289_io_x1 = r_766; // @[MUL.scala 103:13]
  assign m_289_io_x2 = r_767; // @[MUL.scala 104:13]
  assign m_289_io_x3 = r_768; // @[MUL.scala 105:13]
  assign m_290_io_x1 = r_769; // @[MUL.scala 103:13]
  assign m_290_io_x2 = r_770; // @[MUL.scala 104:13]
  assign m_290_io_x3 = r_771; // @[MUL.scala 105:13]
  assign m_291_io_x1 = r_772; // @[MUL.scala 103:13]
  assign m_291_io_x2 = r_773; // @[MUL.scala 104:13]
  assign m_291_io_x3 = r_774; // @[MUL.scala 105:13]
  assign m_292_io_x1 = r_775; // @[MUL.scala 103:13]
  assign m_292_io_x2 = r_776; // @[MUL.scala 104:13]
  assign m_292_io_x3 = r_777; // @[MUL.scala 105:13]
  assign m_293_io_x1 = r_778; // @[MUL.scala 103:13]
  assign m_293_io_x2 = r_779; // @[MUL.scala 104:13]
  assign m_293_io_x3 = r_780; // @[MUL.scala 105:13]
  assign m_294_io_x1 = r_782; // @[MUL.scala 103:13]
  assign m_294_io_x2 = r_783; // @[MUL.scala 104:13]
  assign m_294_io_x3 = r_784; // @[MUL.scala 105:13]
  assign m_295_io_x1 = r_785; // @[MUL.scala 103:13]
  assign m_295_io_x2 = r_786; // @[MUL.scala 104:13]
  assign m_295_io_x3 = r_787; // @[MUL.scala 105:13]
  assign m_296_io_x1 = r_788; // @[MUL.scala 103:13]
  assign m_296_io_x2 = r_789; // @[MUL.scala 104:13]
  assign m_296_io_x3 = r_790; // @[MUL.scala 105:13]
  assign m_297_io_x1 = r_791; // @[MUL.scala 103:13]
  assign m_297_io_x2 = r_792; // @[MUL.scala 104:13]
  assign m_297_io_x3 = r_793; // @[MUL.scala 105:13]
  assign m_298_io_x1 = r_794; // @[MUL.scala 103:13]
  assign m_298_io_x2 = r_795; // @[MUL.scala 104:13]
  assign m_298_io_x3 = r_796; // @[MUL.scala 105:13]
  assign m_299_io_x1 = r_797; // @[MUL.scala 103:13]
  assign m_299_io_x2 = r_798; // @[MUL.scala 104:13]
  assign m_299_io_x3 = r_799; // @[MUL.scala 105:13]
  assign m_300_io_x1 = r_800; // @[MUL.scala 103:13]
  assign m_300_io_x2 = r_801; // @[MUL.scala 104:13]
  assign m_300_io_x3 = r_802; // @[MUL.scala 105:13]
  assign m_301_io_x1 = r_803; // @[MUL.scala 103:13]
  assign m_301_io_x2 = r_804; // @[MUL.scala 104:13]
  assign m_301_io_x3 = r_805; // @[MUL.scala 105:13]
  assign m_302_io_x1 = r_806; // @[MUL.scala 103:13]
  assign m_302_io_x2 = r_807; // @[MUL.scala 104:13]
  assign m_302_io_x3 = r_808; // @[MUL.scala 105:13]
  assign m_303_io_x1 = r_810; // @[MUL.scala 103:13]
  assign m_303_io_x2 = r_811; // @[MUL.scala 104:13]
  assign m_303_io_x3 = r_812; // @[MUL.scala 105:13]
  assign m_304_io_x1 = r_813; // @[MUL.scala 103:13]
  assign m_304_io_x2 = r_814; // @[MUL.scala 104:13]
  assign m_304_io_x3 = r_815; // @[MUL.scala 105:13]
  assign m_305_io_x1 = r_816; // @[MUL.scala 103:13]
  assign m_305_io_x2 = r_817; // @[MUL.scala 104:13]
  assign m_305_io_x3 = r_818; // @[MUL.scala 105:13]
  assign m_306_io_x1 = r_819; // @[MUL.scala 103:13]
  assign m_306_io_x2 = r_820; // @[MUL.scala 104:13]
  assign m_306_io_x3 = r_821; // @[MUL.scala 105:13]
  assign m_307_io_x1 = r_822; // @[MUL.scala 103:13]
  assign m_307_io_x2 = r_823; // @[MUL.scala 104:13]
  assign m_307_io_x3 = r_824; // @[MUL.scala 105:13]
  assign m_308_io_x1 = r_825; // @[MUL.scala 103:13]
  assign m_308_io_x2 = r_826; // @[MUL.scala 104:13]
  assign m_308_io_x3 = r_827; // @[MUL.scala 105:13]
  assign m_309_io_x1 = r_828; // @[MUL.scala 103:13]
  assign m_309_io_x2 = r_829; // @[MUL.scala 104:13]
  assign m_309_io_x3 = r_830; // @[MUL.scala 105:13]
  assign m_310_io_x1 = r_831; // @[MUL.scala 103:13]
  assign m_310_io_x2 = r_832; // @[MUL.scala 104:13]
  assign m_310_io_x3 = r_833; // @[MUL.scala 105:13]
  assign m_311_io_x1 = r_834; // @[MUL.scala 103:13]
  assign m_311_io_x2 = r_835; // @[MUL.scala 104:13]
  assign m_311_io_x3 = r_836; // @[MUL.scala 105:13]
  assign m_312_io_in_0 = r_837; // @[MUL.scala 125:16]
  assign m_312_io_in_1 = r_838; // @[MUL.scala 126:16]
  assign m_313_io_x1 = r_839; // @[MUL.scala 103:13]
  assign m_313_io_x2 = r_840; // @[MUL.scala 104:13]
  assign m_313_io_x3 = r_841; // @[MUL.scala 105:13]
  assign m_314_io_x1 = r_842; // @[MUL.scala 103:13]
  assign m_314_io_x2 = r_843; // @[MUL.scala 104:13]
  assign m_314_io_x3 = r_844; // @[MUL.scala 105:13]
  assign m_315_io_x1 = r_845; // @[MUL.scala 103:13]
  assign m_315_io_x2 = r_846; // @[MUL.scala 104:13]
  assign m_315_io_x3 = r_847; // @[MUL.scala 105:13]
  assign m_316_io_x1 = r_848; // @[MUL.scala 103:13]
  assign m_316_io_x2 = r_849; // @[MUL.scala 104:13]
  assign m_316_io_x3 = r_850; // @[MUL.scala 105:13]
  assign m_317_io_x1 = r_851; // @[MUL.scala 103:13]
  assign m_317_io_x2 = r_852; // @[MUL.scala 104:13]
  assign m_317_io_x3 = r_853; // @[MUL.scala 105:13]
  assign m_318_io_x1 = r_854; // @[MUL.scala 103:13]
  assign m_318_io_x2 = r_855; // @[MUL.scala 104:13]
  assign m_318_io_x3 = r_856; // @[MUL.scala 105:13]
  assign m_319_io_x1 = r_857; // @[MUL.scala 103:13]
  assign m_319_io_x2 = r_858; // @[MUL.scala 104:13]
  assign m_319_io_x3 = r_859; // @[MUL.scala 105:13]
  assign m_320_io_x1 = r_860; // @[MUL.scala 103:13]
  assign m_320_io_x2 = r_861; // @[MUL.scala 104:13]
  assign m_320_io_x3 = r_862; // @[MUL.scala 105:13]
  assign m_321_io_x1 = r_863; // @[MUL.scala 103:13]
  assign m_321_io_x2 = r_864; // @[MUL.scala 104:13]
  assign m_321_io_x3 = r_865; // @[MUL.scala 105:13]
  assign m_322_io_in_0 = r_866; // @[MUL.scala 125:16]
  assign m_322_io_in_1 = r_867; // @[MUL.scala 126:16]
  assign m_323_io_x1 = r_868; // @[MUL.scala 103:13]
  assign m_323_io_x2 = r_869; // @[MUL.scala 104:13]
  assign m_323_io_x3 = r_870; // @[MUL.scala 105:13]
  assign m_324_io_x1 = r_871; // @[MUL.scala 103:13]
  assign m_324_io_x2 = r_872; // @[MUL.scala 104:13]
  assign m_324_io_x3 = r_873; // @[MUL.scala 105:13]
  assign m_325_io_x1 = r_874; // @[MUL.scala 103:13]
  assign m_325_io_x2 = r_875; // @[MUL.scala 104:13]
  assign m_325_io_x3 = r_876; // @[MUL.scala 105:13]
  assign m_326_io_x1 = r_877; // @[MUL.scala 103:13]
  assign m_326_io_x2 = r_878; // @[MUL.scala 104:13]
  assign m_326_io_x3 = r_879; // @[MUL.scala 105:13]
  assign m_327_io_x1 = r_880; // @[MUL.scala 103:13]
  assign m_327_io_x2 = r_881; // @[MUL.scala 104:13]
  assign m_327_io_x3 = r_882; // @[MUL.scala 105:13]
  assign m_328_io_x1 = r_883; // @[MUL.scala 103:13]
  assign m_328_io_x2 = r_884; // @[MUL.scala 104:13]
  assign m_328_io_x3 = r_885; // @[MUL.scala 105:13]
  assign m_329_io_x1 = r_886; // @[MUL.scala 103:13]
  assign m_329_io_x2 = r_887; // @[MUL.scala 104:13]
  assign m_329_io_x3 = r_888; // @[MUL.scala 105:13]
  assign m_330_io_x1 = r_889; // @[MUL.scala 103:13]
  assign m_330_io_x2 = r_890; // @[MUL.scala 104:13]
  assign m_330_io_x3 = r_891; // @[MUL.scala 105:13]
  assign m_331_io_x1 = r_892; // @[MUL.scala 103:13]
  assign m_331_io_x2 = r_893; // @[MUL.scala 104:13]
  assign m_331_io_x3 = r_894; // @[MUL.scala 105:13]
  assign m_332_io_x1 = r_895; // @[MUL.scala 103:13]
  assign m_332_io_x2 = r_896; // @[MUL.scala 104:13]
  assign m_332_io_x3 = r_897; // @[MUL.scala 105:13]
  assign m_333_io_x1 = r_898; // @[MUL.scala 103:13]
  assign m_333_io_x2 = r_899; // @[MUL.scala 104:13]
  assign m_333_io_x3 = r_900; // @[MUL.scala 105:13]
  assign m_334_io_x1 = r_901; // @[MUL.scala 103:13]
  assign m_334_io_x2 = r_902; // @[MUL.scala 104:13]
  assign m_334_io_x3 = r_903; // @[MUL.scala 105:13]
  assign m_335_io_x1 = r_904; // @[MUL.scala 103:13]
  assign m_335_io_x2 = r_905; // @[MUL.scala 104:13]
  assign m_335_io_x3 = r_906; // @[MUL.scala 105:13]
  assign m_336_io_x1 = r_907; // @[MUL.scala 103:13]
  assign m_336_io_x2 = r_908; // @[MUL.scala 104:13]
  assign m_336_io_x3 = r_909; // @[MUL.scala 105:13]
  assign m_337_io_x1 = r_910; // @[MUL.scala 103:13]
  assign m_337_io_x2 = r_911; // @[MUL.scala 104:13]
  assign m_337_io_x3 = r_912; // @[MUL.scala 105:13]
  assign m_338_io_x1 = r_913; // @[MUL.scala 103:13]
  assign m_338_io_x2 = r_914; // @[MUL.scala 104:13]
  assign m_338_io_x3 = r_915; // @[MUL.scala 105:13]
  assign m_339_io_x1 = r_916; // @[MUL.scala 103:13]
  assign m_339_io_x2 = r_917; // @[MUL.scala 104:13]
  assign m_339_io_x3 = r_918; // @[MUL.scala 105:13]
  assign m_340_io_x1 = r_919; // @[MUL.scala 103:13]
  assign m_340_io_x2 = r_920; // @[MUL.scala 104:13]
  assign m_340_io_x3 = r_921; // @[MUL.scala 105:13]
  assign m_341_io_x1 = r_922; // @[MUL.scala 103:13]
  assign m_341_io_x2 = r_923; // @[MUL.scala 104:13]
  assign m_341_io_x3 = r_924; // @[MUL.scala 105:13]
  assign m_342_io_x1 = r_925; // @[MUL.scala 103:13]
  assign m_342_io_x2 = r_926; // @[MUL.scala 104:13]
  assign m_342_io_x3 = r_927; // @[MUL.scala 105:13]
  assign m_343_io_x1 = r_928; // @[MUL.scala 103:13]
  assign m_343_io_x2 = r_929; // @[MUL.scala 104:13]
  assign m_343_io_x3 = r_930; // @[MUL.scala 105:13]
  assign m_344_io_x1 = r_931; // @[MUL.scala 103:13]
  assign m_344_io_x2 = r_932; // @[MUL.scala 104:13]
  assign m_344_io_x3 = r_933; // @[MUL.scala 105:13]
  assign m_345_io_x1 = r_934; // @[MUL.scala 103:13]
  assign m_345_io_x2 = r_935; // @[MUL.scala 104:13]
  assign m_345_io_x3 = r_936; // @[MUL.scala 105:13]
  assign m_346_io_x1 = r_937; // @[MUL.scala 103:13]
  assign m_346_io_x2 = r_938; // @[MUL.scala 104:13]
  assign m_346_io_x3 = r_939; // @[MUL.scala 105:13]
  assign m_347_io_x1 = r_940; // @[MUL.scala 103:13]
  assign m_347_io_x2 = r_941; // @[MUL.scala 104:13]
  assign m_347_io_x3 = r_942; // @[MUL.scala 105:13]
  assign m_348_io_x1 = r_943; // @[MUL.scala 103:13]
  assign m_348_io_x2 = r_944; // @[MUL.scala 104:13]
  assign m_348_io_x3 = r_945; // @[MUL.scala 105:13]
  assign m_349_io_x1 = r_946; // @[MUL.scala 103:13]
  assign m_349_io_x2 = r_947; // @[MUL.scala 104:13]
  assign m_349_io_x3 = r_948; // @[MUL.scala 105:13]
  assign m_350_io_x1 = r_949; // @[MUL.scala 103:13]
  assign m_350_io_x2 = r_950; // @[MUL.scala 104:13]
  assign m_350_io_x3 = r_951; // @[MUL.scala 105:13]
  assign m_351_io_x1 = r_952; // @[MUL.scala 103:13]
  assign m_351_io_x2 = r_953; // @[MUL.scala 104:13]
  assign m_351_io_x3 = r_954; // @[MUL.scala 105:13]
  assign m_352_io_x1 = r_955; // @[MUL.scala 103:13]
  assign m_352_io_x2 = r_956; // @[MUL.scala 104:13]
  assign m_352_io_x3 = r_957; // @[MUL.scala 105:13]
  assign m_353_io_x1 = r_959; // @[MUL.scala 103:13]
  assign m_353_io_x2 = r_960; // @[MUL.scala 104:13]
  assign m_353_io_x3 = r_961; // @[MUL.scala 105:13]
  assign m_354_io_x1 = r_962; // @[MUL.scala 103:13]
  assign m_354_io_x2 = r_963; // @[MUL.scala 104:13]
  assign m_354_io_x3 = r_964; // @[MUL.scala 105:13]
  assign m_355_io_x1 = r_965; // @[MUL.scala 103:13]
  assign m_355_io_x2 = r_966; // @[MUL.scala 104:13]
  assign m_355_io_x3 = r_967; // @[MUL.scala 105:13]
  assign m_356_io_x1 = r_968; // @[MUL.scala 103:13]
  assign m_356_io_x2 = r_969; // @[MUL.scala 104:13]
  assign m_356_io_x3 = r_970; // @[MUL.scala 105:13]
  assign m_357_io_x1 = r_971; // @[MUL.scala 103:13]
  assign m_357_io_x2 = r_972; // @[MUL.scala 104:13]
  assign m_357_io_x3 = r_973; // @[MUL.scala 105:13]
  assign m_358_io_x1 = r_974; // @[MUL.scala 103:13]
  assign m_358_io_x2 = r_975; // @[MUL.scala 104:13]
  assign m_358_io_x3 = r_976; // @[MUL.scala 105:13]
  assign m_359_io_x1 = r_977; // @[MUL.scala 103:13]
  assign m_359_io_x2 = r_978; // @[MUL.scala 104:13]
  assign m_359_io_x3 = r_979; // @[MUL.scala 105:13]
  assign m_360_io_x1 = r_980; // @[MUL.scala 103:13]
  assign m_360_io_x2 = r_981; // @[MUL.scala 104:13]
  assign m_360_io_x3 = r_982; // @[MUL.scala 105:13]
  assign m_361_io_x1 = r_983; // @[MUL.scala 103:13]
  assign m_361_io_x2 = r_984; // @[MUL.scala 104:13]
  assign m_361_io_x3 = r_985; // @[MUL.scala 105:13]
  assign m_362_io_x1 = r_986; // @[MUL.scala 103:13]
  assign m_362_io_x2 = r_987; // @[MUL.scala 104:13]
  assign m_362_io_x3 = r_988; // @[MUL.scala 105:13]
  assign m_363_io_x1 = r_990; // @[MUL.scala 103:13]
  assign m_363_io_x2 = r_991; // @[MUL.scala 104:13]
  assign m_363_io_x3 = r_992; // @[MUL.scala 105:13]
  assign m_364_io_x1 = r_993; // @[MUL.scala 103:13]
  assign m_364_io_x2 = r_994; // @[MUL.scala 104:13]
  assign m_364_io_x3 = r_995; // @[MUL.scala 105:13]
  assign m_365_io_x1 = r_996; // @[MUL.scala 103:13]
  assign m_365_io_x2 = r_997; // @[MUL.scala 104:13]
  assign m_365_io_x3 = r_998; // @[MUL.scala 105:13]
  assign m_366_io_x1 = r_999; // @[MUL.scala 103:13]
  assign m_366_io_x2 = r_1000; // @[MUL.scala 104:13]
  assign m_366_io_x3 = r_1001; // @[MUL.scala 105:13]
  assign m_367_io_x1 = r_1002; // @[MUL.scala 103:13]
  assign m_367_io_x2 = r_1003; // @[MUL.scala 104:13]
  assign m_367_io_x3 = r_1004; // @[MUL.scala 105:13]
  assign m_368_io_x1 = r_1005; // @[MUL.scala 103:13]
  assign m_368_io_x2 = r_1006; // @[MUL.scala 104:13]
  assign m_368_io_x3 = r_1007; // @[MUL.scala 105:13]
  assign m_369_io_x1 = r_1008; // @[MUL.scala 103:13]
  assign m_369_io_x2 = r_1009; // @[MUL.scala 104:13]
  assign m_369_io_x3 = r_1010; // @[MUL.scala 105:13]
  assign m_370_io_x1 = r_1011; // @[MUL.scala 103:13]
  assign m_370_io_x2 = r_1012; // @[MUL.scala 104:13]
  assign m_370_io_x3 = r_1013; // @[MUL.scala 105:13]
  assign m_371_io_x1 = r_1014; // @[MUL.scala 103:13]
  assign m_371_io_x2 = r_1015; // @[MUL.scala 104:13]
  assign m_371_io_x3 = r_1016; // @[MUL.scala 105:13]
  assign m_372_io_x1 = r_1017; // @[MUL.scala 103:13]
  assign m_372_io_x2 = r_1018; // @[MUL.scala 104:13]
  assign m_372_io_x3 = r_1019; // @[MUL.scala 105:13]
  assign m_373_io_in_0 = r_1020; // @[MUL.scala 125:16]
  assign m_373_io_in_1 = r_1021; // @[MUL.scala 126:16]
  assign m_374_io_x1 = r_1022; // @[MUL.scala 103:13]
  assign m_374_io_x2 = r_1023; // @[MUL.scala 104:13]
  assign m_374_io_x3 = r_1024; // @[MUL.scala 105:13]
  assign m_375_io_x1 = r_1025; // @[MUL.scala 103:13]
  assign m_375_io_x2 = r_1026; // @[MUL.scala 104:13]
  assign m_375_io_x3 = r_1027; // @[MUL.scala 105:13]
  assign m_376_io_x1 = r_1028; // @[MUL.scala 103:13]
  assign m_376_io_x2 = r_1029; // @[MUL.scala 104:13]
  assign m_376_io_x3 = r_1030; // @[MUL.scala 105:13]
  assign m_377_io_x1 = r_1031; // @[MUL.scala 103:13]
  assign m_377_io_x2 = r_1032; // @[MUL.scala 104:13]
  assign m_377_io_x3 = r_1033; // @[MUL.scala 105:13]
  assign m_378_io_x1 = r_1034; // @[MUL.scala 103:13]
  assign m_378_io_x2 = r_1035; // @[MUL.scala 104:13]
  assign m_378_io_x3 = r_1036; // @[MUL.scala 105:13]
  assign m_379_io_x1 = r_1037; // @[MUL.scala 103:13]
  assign m_379_io_x2 = r_1038; // @[MUL.scala 104:13]
  assign m_379_io_x3 = r_1039; // @[MUL.scala 105:13]
  assign m_380_io_x1 = r_1040; // @[MUL.scala 103:13]
  assign m_380_io_x2 = r_1041; // @[MUL.scala 104:13]
  assign m_380_io_x3 = r_1042; // @[MUL.scala 105:13]
  assign m_381_io_x1 = r_1043; // @[MUL.scala 103:13]
  assign m_381_io_x2 = r_1044; // @[MUL.scala 104:13]
  assign m_381_io_x3 = r_1045; // @[MUL.scala 105:13]
  assign m_382_io_x1 = r_1046; // @[MUL.scala 103:13]
  assign m_382_io_x2 = r_1047; // @[MUL.scala 104:13]
  assign m_382_io_x3 = r_1048; // @[MUL.scala 105:13]
  assign m_383_io_x1 = r_1049; // @[MUL.scala 103:13]
  assign m_383_io_x2 = r_1050; // @[MUL.scala 104:13]
  assign m_383_io_x3 = r_1051; // @[MUL.scala 105:13]
  assign m_384_io_in_0 = r_1052; // @[MUL.scala 125:16]
  assign m_384_io_in_1 = r_1053; // @[MUL.scala 126:16]
  assign m_385_io_x1 = r_1054; // @[MUL.scala 103:13]
  assign m_385_io_x2 = r_1055; // @[MUL.scala 104:13]
  assign m_385_io_x3 = r_1056; // @[MUL.scala 105:13]
  assign m_386_io_x1 = r_1057; // @[MUL.scala 103:13]
  assign m_386_io_x2 = r_1058; // @[MUL.scala 104:13]
  assign m_386_io_x3 = r_1059; // @[MUL.scala 105:13]
  assign m_387_io_x1 = r_1060; // @[MUL.scala 103:13]
  assign m_387_io_x2 = r_1061; // @[MUL.scala 104:13]
  assign m_387_io_x3 = r_1062; // @[MUL.scala 105:13]
  assign m_388_io_x1 = r_1063; // @[MUL.scala 103:13]
  assign m_388_io_x2 = r_1064; // @[MUL.scala 104:13]
  assign m_388_io_x3 = r_1065; // @[MUL.scala 105:13]
  assign m_389_io_x1 = r_1066; // @[MUL.scala 103:13]
  assign m_389_io_x2 = r_1067; // @[MUL.scala 104:13]
  assign m_389_io_x3 = r_1068; // @[MUL.scala 105:13]
  assign m_390_io_x1 = r_1069; // @[MUL.scala 103:13]
  assign m_390_io_x2 = r_1070; // @[MUL.scala 104:13]
  assign m_390_io_x3 = r_1071; // @[MUL.scala 105:13]
  assign m_391_io_x1 = r_1072; // @[MUL.scala 103:13]
  assign m_391_io_x2 = r_1073; // @[MUL.scala 104:13]
  assign m_391_io_x3 = r_1074; // @[MUL.scala 105:13]
  assign m_392_io_x1 = r_1075; // @[MUL.scala 103:13]
  assign m_392_io_x2 = r_1076; // @[MUL.scala 104:13]
  assign m_392_io_x3 = r_1077; // @[MUL.scala 105:13]
  assign m_393_io_x1 = r_1078; // @[MUL.scala 103:13]
  assign m_393_io_x2 = r_1079; // @[MUL.scala 104:13]
  assign m_393_io_x3 = r_1080; // @[MUL.scala 105:13]
  assign m_394_io_x1 = r_1081; // @[MUL.scala 103:13]
  assign m_394_io_x2 = r_1082; // @[MUL.scala 104:13]
  assign m_394_io_x3 = r_1083; // @[MUL.scala 105:13]
  assign m_395_io_x1 = r_1084; // @[MUL.scala 103:13]
  assign m_395_io_x2 = r_1085; // @[MUL.scala 104:13]
  assign m_395_io_x3 = r_1086; // @[MUL.scala 105:13]
  assign m_396_io_x1 = r_1087; // @[MUL.scala 103:13]
  assign m_396_io_x2 = r_1088; // @[MUL.scala 104:13]
  assign m_396_io_x3 = r_1089; // @[MUL.scala 105:13]
  assign m_397_io_x1 = r_1090; // @[MUL.scala 103:13]
  assign m_397_io_x2 = r_1091; // @[MUL.scala 104:13]
  assign m_397_io_x3 = r_1092; // @[MUL.scala 105:13]
  assign m_398_io_x1 = r_1093; // @[MUL.scala 103:13]
  assign m_398_io_x2 = r_1094; // @[MUL.scala 104:13]
  assign m_398_io_x3 = r_1095; // @[MUL.scala 105:13]
  assign m_399_io_x1 = r_1096; // @[MUL.scala 103:13]
  assign m_399_io_x2 = r_1097; // @[MUL.scala 104:13]
  assign m_399_io_x3 = r_1098; // @[MUL.scala 105:13]
  assign m_400_io_x1 = r_1099; // @[MUL.scala 103:13]
  assign m_400_io_x2 = r_1100; // @[MUL.scala 104:13]
  assign m_400_io_x3 = r_1101; // @[MUL.scala 105:13]
  assign m_401_io_x1 = r_1102; // @[MUL.scala 103:13]
  assign m_401_io_x2 = r_1103; // @[MUL.scala 104:13]
  assign m_401_io_x3 = r_1104; // @[MUL.scala 105:13]
  assign m_402_io_x1 = r_1105; // @[MUL.scala 103:13]
  assign m_402_io_x2 = r_1106; // @[MUL.scala 104:13]
  assign m_402_io_x3 = r_1107; // @[MUL.scala 105:13]
  assign m_403_io_x1 = r_1108; // @[MUL.scala 103:13]
  assign m_403_io_x2 = r_1109; // @[MUL.scala 104:13]
  assign m_403_io_x3 = r_1110; // @[MUL.scala 105:13]
  assign m_404_io_x1 = r_1111; // @[MUL.scala 103:13]
  assign m_404_io_x2 = r_1112; // @[MUL.scala 104:13]
  assign m_404_io_x3 = r_1113; // @[MUL.scala 105:13]
  assign m_405_io_x1 = r_1114; // @[MUL.scala 103:13]
  assign m_405_io_x2 = r_1115; // @[MUL.scala 104:13]
  assign m_405_io_x3 = r_1116; // @[MUL.scala 105:13]
  assign m_406_io_x1 = r_1117; // @[MUL.scala 103:13]
  assign m_406_io_x2 = r_1118; // @[MUL.scala 104:13]
  assign m_406_io_x3 = r_1119; // @[MUL.scala 105:13]
  assign m_407_io_x1 = r_1120; // @[MUL.scala 103:13]
  assign m_407_io_x2 = r_1121; // @[MUL.scala 104:13]
  assign m_407_io_x3 = r_1122; // @[MUL.scala 105:13]
  assign m_408_io_x1 = r_1123; // @[MUL.scala 103:13]
  assign m_408_io_x2 = r_1124; // @[MUL.scala 104:13]
  assign m_408_io_x3 = r_1125; // @[MUL.scala 105:13]
  assign m_409_io_x1 = r_1126; // @[MUL.scala 103:13]
  assign m_409_io_x2 = r_1127; // @[MUL.scala 104:13]
  assign m_409_io_x3 = r_1128; // @[MUL.scala 105:13]
  assign m_410_io_x1 = r_1129; // @[MUL.scala 103:13]
  assign m_410_io_x2 = r_1130; // @[MUL.scala 104:13]
  assign m_410_io_x3 = r_1131; // @[MUL.scala 105:13]
  assign m_411_io_x1 = r_1132; // @[MUL.scala 103:13]
  assign m_411_io_x2 = r_1133; // @[MUL.scala 104:13]
  assign m_411_io_x3 = r_1134; // @[MUL.scala 105:13]
  assign m_412_io_x1 = r_1135; // @[MUL.scala 103:13]
  assign m_412_io_x2 = r_1136; // @[MUL.scala 104:13]
  assign m_412_io_x3 = r_1137; // @[MUL.scala 105:13]
  assign m_413_io_x1 = r_1138; // @[MUL.scala 103:13]
  assign m_413_io_x2 = r_1139; // @[MUL.scala 104:13]
  assign m_413_io_x3 = r_1140; // @[MUL.scala 105:13]
  assign m_414_io_x1 = r_1141; // @[MUL.scala 103:13]
  assign m_414_io_x2 = r_1142; // @[MUL.scala 104:13]
  assign m_414_io_x3 = r_1143; // @[MUL.scala 105:13]
  assign m_415_io_x1 = r_1144; // @[MUL.scala 103:13]
  assign m_415_io_x2 = r_1145; // @[MUL.scala 104:13]
  assign m_415_io_x3 = r_1146; // @[MUL.scala 105:13]
  assign m_416_io_x1 = r_1147; // @[MUL.scala 103:13]
  assign m_416_io_x2 = r_1148; // @[MUL.scala 104:13]
  assign m_416_io_x3 = r_1149; // @[MUL.scala 105:13]
  assign m_417_io_x1 = r_1150; // @[MUL.scala 103:13]
  assign m_417_io_x2 = r_1151; // @[MUL.scala 104:13]
  assign m_417_io_x3 = r_1152; // @[MUL.scala 105:13]
  assign m_418_io_x1 = r_1153; // @[MUL.scala 103:13]
  assign m_418_io_x2 = r_1154; // @[MUL.scala 104:13]
  assign m_418_io_x3 = r_1155; // @[MUL.scala 105:13]
  assign m_419_io_x1 = r_1156; // @[MUL.scala 103:13]
  assign m_419_io_x2 = r_1157; // @[MUL.scala 104:13]
  assign m_419_io_x3 = r_1158; // @[MUL.scala 105:13]
  assign m_420_io_x1 = r_1159; // @[MUL.scala 103:13]
  assign m_420_io_x2 = r_1160; // @[MUL.scala 104:13]
  assign m_420_io_x3 = r_1161; // @[MUL.scala 105:13]
  assign m_421_io_x1 = r_1162; // @[MUL.scala 103:13]
  assign m_421_io_x2 = r_1163; // @[MUL.scala 104:13]
  assign m_421_io_x3 = r_1164; // @[MUL.scala 105:13]
  assign m_422_io_x1 = r_1165; // @[MUL.scala 103:13]
  assign m_422_io_x2 = r_1166; // @[MUL.scala 104:13]
  assign m_422_io_x3 = r_1167; // @[MUL.scala 105:13]
  assign m_423_io_x1 = r_1168; // @[MUL.scala 103:13]
  assign m_423_io_x2 = r_1169; // @[MUL.scala 104:13]
  assign m_423_io_x3 = r_1170; // @[MUL.scala 105:13]
  assign m_424_io_x1 = r_1171; // @[MUL.scala 103:13]
  assign m_424_io_x2 = r_1172; // @[MUL.scala 104:13]
  assign m_424_io_x3 = r_1173; // @[MUL.scala 105:13]
  assign m_425_io_x1 = r_1174; // @[MUL.scala 103:13]
  assign m_425_io_x2 = r_1175; // @[MUL.scala 104:13]
  assign m_425_io_x3 = r_1176; // @[MUL.scala 105:13]
  assign m_426_io_x1 = r_1177; // @[MUL.scala 103:13]
  assign m_426_io_x2 = r_1178; // @[MUL.scala 104:13]
  assign m_426_io_x3 = r_1179; // @[MUL.scala 105:13]
  assign m_427_io_x1 = r_1180; // @[MUL.scala 103:13]
  assign m_427_io_x2 = r_1181; // @[MUL.scala 104:13]
  assign m_427_io_x3 = r_1182; // @[MUL.scala 105:13]
  assign m_428_io_x1 = r_1183; // @[MUL.scala 103:13]
  assign m_428_io_x2 = r_1184; // @[MUL.scala 104:13]
  assign m_428_io_x3 = r_1185; // @[MUL.scala 105:13]
  assign m_429_io_x1 = r_1186; // @[MUL.scala 103:13]
  assign m_429_io_x2 = r_1187; // @[MUL.scala 104:13]
  assign m_429_io_x3 = r_1188; // @[MUL.scala 105:13]
  assign m_430_io_x1 = r_1189; // @[MUL.scala 103:13]
  assign m_430_io_x2 = r_1190; // @[MUL.scala 104:13]
  assign m_430_io_x3 = r_1191; // @[MUL.scala 105:13]
  assign m_431_io_x1 = r_1192; // @[MUL.scala 103:13]
  assign m_431_io_x2 = r_1193; // @[MUL.scala 104:13]
  assign m_431_io_x3 = r_1194; // @[MUL.scala 105:13]
  assign m_432_io_x1 = r_1195; // @[MUL.scala 103:13]
  assign m_432_io_x2 = r_1196; // @[MUL.scala 104:13]
  assign m_432_io_x3 = r_1197; // @[MUL.scala 105:13]
  assign m_433_io_x1 = r_1198; // @[MUL.scala 103:13]
  assign m_433_io_x2 = r_1199; // @[MUL.scala 104:13]
  assign m_433_io_x3 = r_1200; // @[MUL.scala 105:13]
  assign m_434_io_x1 = r_1201; // @[MUL.scala 103:13]
  assign m_434_io_x2 = r_1202; // @[MUL.scala 104:13]
  assign m_434_io_x3 = r_1203; // @[MUL.scala 105:13]
  assign m_435_io_x1 = r_1204; // @[MUL.scala 103:13]
  assign m_435_io_x2 = r_1205; // @[MUL.scala 104:13]
  assign m_435_io_x3 = r_1206; // @[MUL.scala 105:13]
  assign m_436_io_x1 = r_1207; // @[MUL.scala 103:13]
  assign m_436_io_x2 = r_1208; // @[MUL.scala 104:13]
  assign m_436_io_x3 = r_1209; // @[MUL.scala 105:13]
  assign m_437_io_x1 = r_1210; // @[MUL.scala 103:13]
  assign m_437_io_x2 = r_1211; // @[MUL.scala 104:13]
  assign m_437_io_x3 = r_1212; // @[MUL.scala 105:13]
  assign m_438_io_x1 = r_1213; // @[MUL.scala 103:13]
  assign m_438_io_x2 = r_1214; // @[MUL.scala 104:13]
  assign m_438_io_x3 = r_1215; // @[MUL.scala 105:13]
  assign m_439_io_x1 = r_1216; // @[MUL.scala 103:13]
  assign m_439_io_x2 = r_1217; // @[MUL.scala 104:13]
  assign m_439_io_x3 = r_1218; // @[MUL.scala 105:13]
  assign m_440_io_x1 = r_1219; // @[MUL.scala 103:13]
  assign m_440_io_x2 = r_1220; // @[MUL.scala 104:13]
  assign m_440_io_x3 = r_1221; // @[MUL.scala 105:13]
  assign m_441_io_x1 = r_1222; // @[MUL.scala 103:13]
  assign m_441_io_x2 = r_1223; // @[MUL.scala 104:13]
  assign m_441_io_x3 = r_1224; // @[MUL.scala 105:13]
  assign m_442_io_x1 = r_1225; // @[MUL.scala 103:13]
  assign m_442_io_x2 = r_1226; // @[MUL.scala 104:13]
  assign m_442_io_x3 = r_1227; // @[MUL.scala 105:13]
  assign m_443_io_x1 = r_1228; // @[MUL.scala 103:13]
  assign m_443_io_x2 = r_1229; // @[MUL.scala 104:13]
  assign m_443_io_x3 = r_1230; // @[MUL.scala 105:13]
  assign m_444_io_x1 = r_1231; // @[MUL.scala 103:13]
  assign m_444_io_x2 = r_1232; // @[MUL.scala 104:13]
  assign m_444_io_x3 = r_1233; // @[MUL.scala 105:13]
  assign m_445_io_x1 = r_1234; // @[MUL.scala 103:13]
  assign m_445_io_x2 = r_1235; // @[MUL.scala 104:13]
  assign m_445_io_x3 = r_1236; // @[MUL.scala 105:13]
  assign m_446_io_x1 = r_1237; // @[MUL.scala 103:13]
  assign m_446_io_x2 = r_1238; // @[MUL.scala 104:13]
  assign m_446_io_x3 = r_1239; // @[MUL.scala 105:13]
  assign m_447_io_x1 = r_1240; // @[MUL.scala 103:13]
  assign m_447_io_x2 = r_1241; // @[MUL.scala 104:13]
  assign m_447_io_x3 = r_1242; // @[MUL.scala 105:13]
  assign m_448_io_x1 = r_1243; // @[MUL.scala 103:13]
  assign m_448_io_x2 = r_1244; // @[MUL.scala 104:13]
  assign m_448_io_x3 = r_1245; // @[MUL.scala 105:13]
  assign m_449_io_x1 = r_1246; // @[MUL.scala 103:13]
  assign m_449_io_x2 = r_1247; // @[MUL.scala 104:13]
  assign m_449_io_x3 = r_1248; // @[MUL.scala 105:13]
  assign m_450_io_x1 = r_1249; // @[MUL.scala 103:13]
  assign m_450_io_x2 = r_1250; // @[MUL.scala 104:13]
  assign m_450_io_x3 = r_1251; // @[MUL.scala 105:13]
  assign m_451_io_x1 = r_1252; // @[MUL.scala 103:13]
  assign m_451_io_x2 = r_1253; // @[MUL.scala 104:13]
  assign m_451_io_x3 = r_1254; // @[MUL.scala 105:13]
  assign m_452_io_x1 = r_1255; // @[MUL.scala 103:13]
  assign m_452_io_x2 = r_1256; // @[MUL.scala 104:13]
  assign m_452_io_x3 = r_1257; // @[MUL.scala 105:13]
  assign m_453_io_x1 = r_1258; // @[MUL.scala 103:13]
  assign m_453_io_x2 = r_1259; // @[MUL.scala 104:13]
  assign m_453_io_x3 = r_1260; // @[MUL.scala 105:13]
  assign m_454_io_x1 = r_1261; // @[MUL.scala 103:13]
  assign m_454_io_x2 = r_1262; // @[MUL.scala 104:13]
  assign m_454_io_x3 = r_1263; // @[MUL.scala 105:13]
  assign m_455_io_x1 = r_1264; // @[MUL.scala 103:13]
  assign m_455_io_x2 = r_1265; // @[MUL.scala 104:13]
  assign m_455_io_x3 = r_1266; // @[MUL.scala 105:13]
  assign m_456_io_x1 = r_1267; // @[MUL.scala 103:13]
  assign m_456_io_x2 = r_1268; // @[MUL.scala 104:13]
  assign m_456_io_x3 = r_1269; // @[MUL.scala 105:13]
  assign m_457_io_x1 = r_1270; // @[MUL.scala 103:13]
  assign m_457_io_x2 = r_1271; // @[MUL.scala 104:13]
  assign m_457_io_x3 = r_1272; // @[MUL.scala 105:13]
  assign m_458_io_x1 = r_1273; // @[MUL.scala 103:13]
  assign m_458_io_x2 = r_1274; // @[MUL.scala 104:13]
  assign m_458_io_x3 = r_1275; // @[MUL.scala 105:13]
  assign m_459_io_x1 = r_1276; // @[MUL.scala 103:13]
  assign m_459_io_x2 = r_1277; // @[MUL.scala 104:13]
  assign m_459_io_x3 = r_1278; // @[MUL.scala 105:13]
  assign m_460_io_x1 = r_1279; // @[MUL.scala 103:13]
  assign m_460_io_x2 = r_1280; // @[MUL.scala 104:13]
  assign m_460_io_x3 = r_1281; // @[MUL.scala 105:13]
  assign m_461_io_x1 = r_1282; // @[MUL.scala 103:13]
  assign m_461_io_x2 = r_1283; // @[MUL.scala 104:13]
  assign m_461_io_x3 = r_1284; // @[MUL.scala 105:13]
  assign m_462_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_462_io_x2 = r_1286; // @[MUL.scala 104:13]
  assign m_462_io_x3 = r_1287; // @[MUL.scala 105:13]
  assign m_463_io_x1 = r_1288; // @[MUL.scala 103:13]
  assign m_463_io_x2 = r_1289; // @[MUL.scala 104:13]
  assign m_463_io_x3 = r_1290; // @[MUL.scala 105:13]
  assign m_464_io_x1 = r_1291; // @[MUL.scala 103:13]
  assign m_464_io_x2 = r_1292; // @[MUL.scala 104:13]
  assign m_464_io_x3 = r_1293; // @[MUL.scala 105:13]
  assign m_465_io_x1 = r_1294; // @[MUL.scala 103:13]
  assign m_465_io_x2 = r_1295; // @[MUL.scala 104:13]
  assign m_465_io_x3 = r_1296; // @[MUL.scala 105:13]
  assign m_466_io_x1 = r_1297; // @[MUL.scala 103:13]
  assign m_466_io_x2 = r_1298; // @[MUL.scala 104:13]
  assign m_466_io_x3 = r_1299; // @[MUL.scala 105:13]
  assign m_467_io_x1 = r_1300; // @[MUL.scala 103:13]
  assign m_467_io_x2 = r_1301; // @[MUL.scala 104:13]
  assign m_467_io_x3 = r_1302; // @[MUL.scala 105:13]
  assign m_468_io_x1 = r_1303; // @[MUL.scala 103:13]
  assign m_468_io_x2 = r_1304; // @[MUL.scala 104:13]
  assign m_468_io_x3 = r_1305; // @[MUL.scala 105:13]
  assign m_469_io_x1 = r_1306; // @[MUL.scala 103:13]
  assign m_469_io_x2 = r_1307; // @[MUL.scala 104:13]
  assign m_469_io_x3 = r_1308; // @[MUL.scala 105:13]
  assign m_470_io_x1 = r_1309; // @[MUL.scala 103:13]
  assign m_470_io_x2 = r_1310; // @[MUL.scala 104:13]
  assign m_470_io_x3 = r_1311; // @[MUL.scala 105:13]
  assign m_471_io_x1 = r_1312; // @[MUL.scala 103:13]
  assign m_471_io_x2 = r_1313; // @[MUL.scala 104:13]
  assign m_471_io_x3 = r_1314; // @[MUL.scala 105:13]
  assign m_472_io_in_0 = r_1315; // @[MUL.scala 125:16]
  assign m_472_io_in_1 = r_1316; // @[MUL.scala 126:16]
  assign m_473_io_x1 = r_1317; // @[MUL.scala 103:13]
  assign m_473_io_x2 = r_1318; // @[MUL.scala 104:13]
  assign m_473_io_x3 = r_1319; // @[MUL.scala 105:13]
  assign m_474_io_x1 = r_1320; // @[MUL.scala 103:13]
  assign m_474_io_x2 = r_1321; // @[MUL.scala 104:13]
  assign m_474_io_x3 = r_1322; // @[MUL.scala 105:13]
  assign m_475_io_x1 = r_1323; // @[MUL.scala 103:13]
  assign m_475_io_x2 = r_1324; // @[MUL.scala 104:13]
  assign m_475_io_x3 = r_1325; // @[MUL.scala 105:13]
  assign m_476_io_x1 = r_1326; // @[MUL.scala 103:13]
  assign m_476_io_x2 = r_1327; // @[MUL.scala 104:13]
  assign m_476_io_x3 = r_1328; // @[MUL.scala 105:13]
  assign m_477_io_x1 = r_1329; // @[MUL.scala 103:13]
  assign m_477_io_x2 = r_1330; // @[MUL.scala 104:13]
  assign m_477_io_x3 = r_1331; // @[MUL.scala 105:13]
  assign m_478_io_x1 = r_1332; // @[MUL.scala 103:13]
  assign m_478_io_x2 = r_1333; // @[MUL.scala 104:13]
  assign m_478_io_x3 = r_1334; // @[MUL.scala 105:13]
  assign m_479_io_x1 = r_1335; // @[MUL.scala 103:13]
  assign m_479_io_x2 = r_1336; // @[MUL.scala 104:13]
  assign m_479_io_x3 = r_1337; // @[MUL.scala 105:13]
  assign m_480_io_x1 = r_1338; // @[MUL.scala 103:13]
  assign m_480_io_x2 = r_1339; // @[MUL.scala 104:13]
  assign m_480_io_x3 = r_1340; // @[MUL.scala 105:13]
  assign m_481_io_x1 = r_1341; // @[MUL.scala 103:13]
  assign m_481_io_x2 = r_1342; // @[MUL.scala 104:13]
  assign m_481_io_x3 = r_1343; // @[MUL.scala 105:13]
  assign m_482_io_x1 = r_1344; // @[MUL.scala 103:13]
  assign m_482_io_x2 = r_1345; // @[MUL.scala 104:13]
  assign m_482_io_x3 = r_1346; // @[MUL.scala 105:13]
  assign m_483_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_483_io_x2 = r_1349; // @[MUL.scala 104:13]
  assign m_483_io_x3 = r_1350; // @[MUL.scala 105:13]
  assign m_484_io_x1 = r_1351; // @[MUL.scala 103:13]
  assign m_484_io_x2 = r_1352; // @[MUL.scala 104:13]
  assign m_484_io_x3 = r_1353; // @[MUL.scala 105:13]
  assign m_485_io_x1 = r_1354; // @[MUL.scala 103:13]
  assign m_485_io_x2 = r_1355; // @[MUL.scala 104:13]
  assign m_485_io_x3 = r_1356; // @[MUL.scala 105:13]
  assign m_486_io_x1 = r_1357; // @[MUL.scala 103:13]
  assign m_486_io_x2 = r_1358; // @[MUL.scala 104:13]
  assign m_486_io_x3 = r_1359; // @[MUL.scala 105:13]
  assign m_487_io_x1 = r_1360; // @[MUL.scala 103:13]
  assign m_487_io_x2 = r_1361; // @[MUL.scala 104:13]
  assign m_487_io_x3 = r_1362; // @[MUL.scala 105:13]
  assign m_488_io_x1 = r_1363; // @[MUL.scala 103:13]
  assign m_488_io_x2 = r_1364; // @[MUL.scala 104:13]
  assign m_488_io_x3 = r_1365; // @[MUL.scala 105:13]
  assign m_489_io_x1 = r_1366; // @[MUL.scala 103:13]
  assign m_489_io_x2 = r_1367; // @[MUL.scala 104:13]
  assign m_489_io_x3 = r_1368; // @[MUL.scala 105:13]
  assign m_490_io_x1 = r_1369; // @[MUL.scala 103:13]
  assign m_490_io_x2 = r_1370; // @[MUL.scala 104:13]
  assign m_490_io_x3 = r_1371; // @[MUL.scala 105:13]
  assign m_491_io_x1 = r_1372; // @[MUL.scala 103:13]
  assign m_491_io_x2 = r_1373; // @[MUL.scala 104:13]
  assign m_491_io_x3 = r_1374; // @[MUL.scala 105:13]
  assign m_492_io_x1 = r_1375; // @[MUL.scala 103:13]
  assign m_492_io_x2 = r_1376; // @[MUL.scala 104:13]
  assign m_492_io_x3 = r_1377; // @[MUL.scala 105:13]
  assign m_493_io_x1 = r_1379; // @[MUL.scala 103:13]
  assign m_493_io_x2 = r_1380; // @[MUL.scala 104:13]
  assign m_493_io_x3 = r_1381; // @[MUL.scala 105:13]
  assign m_494_io_x1 = r_1382; // @[MUL.scala 103:13]
  assign m_494_io_x2 = r_1383; // @[MUL.scala 104:13]
  assign m_494_io_x3 = r_1384; // @[MUL.scala 105:13]
  assign m_495_io_x1 = r_1385; // @[MUL.scala 103:13]
  assign m_495_io_x2 = r_1386; // @[MUL.scala 104:13]
  assign m_495_io_x3 = r_1387; // @[MUL.scala 105:13]
  assign m_496_io_x1 = r_1388; // @[MUL.scala 103:13]
  assign m_496_io_x2 = r_1389; // @[MUL.scala 104:13]
  assign m_496_io_x3 = r_1390; // @[MUL.scala 105:13]
  assign m_497_io_x1 = r_1391; // @[MUL.scala 103:13]
  assign m_497_io_x2 = r_1392; // @[MUL.scala 104:13]
  assign m_497_io_x3 = r_1393; // @[MUL.scala 105:13]
  assign m_498_io_x1 = r_1394; // @[MUL.scala 103:13]
  assign m_498_io_x2 = r_1395; // @[MUL.scala 104:13]
  assign m_498_io_x3 = r_1396; // @[MUL.scala 105:13]
  assign m_499_io_x1 = r_1397; // @[MUL.scala 103:13]
  assign m_499_io_x2 = r_1398; // @[MUL.scala 104:13]
  assign m_499_io_x3 = r_1399; // @[MUL.scala 105:13]
  assign m_500_io_x1 = r_1400; // @[MUL.scala 103:13]
  assign m_500_io_x2 = r_1401; // @[MUL.scala 104:13]
  assign m_500_io_x3 = r_1402; // @[MUL.scala 105:13]
  assign m_501_io_x1 = r_1403; // @[MUL.scala 103:13]
  assign m_501_io_x2 = r_1404; // @[MUL.scala 104:13]
  assign m_501_io_x3 = r_1405; // @[MUL.scala 105:13]
  assign m_502_io_x1 = r_1406; // @[MUL.scala 103:13]
  assign m_502_io_x2 = r_1407; // @[MUL.scala 104:13]
  assign m_502_io_x3 = r_1408; // @[MUL.scala 105:13]
  assign m_503_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_503_io_x2 = r_1410; // @[MUL.scala 104:13]
  assign m_503_io_x3 = r_1411; // @[MUL.scala 105:13]
  assign m_504_io_x1 = r_1412; // @[MUL.scala 103:13]
  assign m_504_io_x2 = r_1413; // @[MUL.scala 104:13]
  assign m_504_io_x3 = r_1414; // @[MUL.scala 105:13]
  assign m_505_io_x1 = r_1415; // @[MUL.scala 103:13]
  assign m_505_io_x2 = r_1416; // @[MUL.scala 104:13]
  assign m_505_io_x3 = r_1417; // @[MUL.scala 105:13]
  assign m_506_io_x1 = r_1418; // @[MUL.scala 103:13]
  assign m_506_io_x2 = r_1419; // @[MUL.scala 104:13]
  assign m_506_io_x3 = r_1420; // @[MUL.scala 105:13]
  assign m_507_io_x1 = r_1421; // @[MUL.scala 103:13]
  assign m_507_io_x2 = r_1422; // @[MUL.scala 104:13]
  assign m_507_io_x3 = r_1423; // @[MUL.scala 105:13]
  assign m_508_io_x1 = r_1424; // @[MUL.scala 103:13]
  assign m_508_io_x2 = r_1425; // @[MUL.scala 104:13]
  assign m_508_io_x3 = r_1426; // @[MUL.scala 105:13]
  assign m_509_io_x1 = r_1427; // @[MUL.scala 103:13]
  assign m_509_io_x2 = r_1428; // @[MUL.scala 104:13]
  assign m_509_io_x3 = r_1429; // @[MUL.scala 105:13]
  assign m_510_io_x1 = r_1430; // @[MUL.scala 103:13]
  assign m_510_io_x2 = r_1431; // @[MUL.scala 104:13]
  assign m_510_io_x3 = r_1432; // @[MUL.scala 105:13]
  assign m_511_io_x1 = r_1433; // @[MUL.scala 103:13]
  assign m_511_io_x2 = r_1434; // @[MUL.scala 104:13]
  assign m_511_io_x3 = r_1435; // @[MUL.scala 105:13]
  assign m_512_io_x1 = r_1436; // @[MUL.scala 103:13]
  assign m_512_io_x2 = r_1437; // @[MUL.scala 104:13]
  assign m_512_io_x3 = r_1438; // @[MUL.scala 105:13]
  assign m_513_io_x1 = r_1439; // @[MUL.scala 103:13]
  assign m_513_io_x2 = r_1440; // @[MUL.scala 104:13]
  assign m_513_io_x3 = r_1441; // @[MUL.scala 105:13]
  assign m_514_io_x1 = r_1442; // @[MUL.scala 103:13]
  assign m_514_io_x2 = r_1443; // @[MUL.scala 104:13]
  assign m_514_io_x3 = r_1444; // @[MUL.scala 105:13]
  assign m_515_io_x1 = r_1445; // @[MUL.scala 103:13]
  assign m_515_io_x2 = r_1446; // @[MUL.scala 104:13]
  assign m_515_io_x3 = r_1447; // @[MUL.scala 105:13]
  assign m_516_io_x1 = r_1448; // @[MUL.scala 103:13]
  assign m_516_io_x2 = r_1449; // @[MUL.scala 104:13]
  assign m_516_io_x3 = r_1450; // @[MUL.scala 105:13]
  assign m_517_io_x1 = r_1451; // @[MUL.scala 103:13]
  assign m_517_io_x2 = r_1452; // @[MUL.scala 104:13]
  assign m_517_io_x3 = r_1453; // @[MUL.scala 105:13]
  assign m_518_io_x1 = r_1454; // @[MUL.scala 103:13]
  assign m_518_io_x2 = r_1455; // @[MUL.scala 104:13]
  assign m_518_io_x3 = r_1456; // @[MUL.scala 105:13]
  assign m_519_io_x1 = r_1457; // @[MUL.scala 103:13]
  assign m_519_io_x2 = r_1458; // @[MUL.scala 104:13]
  assign m_519_io_x3 = r_1459; // @[MUL.scala 105:13]
  assign m_520_io_x1 = r_1460; // @[MUL.scala 103:13]
  assign m_520_io_x2 = r_1461; // @[MUL.scala 104:13]
  assign m_520_io_x3 = r_1462; // @[MUL.scala 105:13]
  assign m_521_io_x1 = r_1463; // @[MUL.scala 103:13]
  assign m_521_io_x2 = r_1464; // @[MUL.scala 104:13]
  assign m_521_io_x3 = r_1465; // @[MUL.scala 105:13]
  assign m_522_io_in_0 = r_1466; // @[MUL.scala 125:16]
  assign m_522_io_in_1 = r_1467; // @[MUL.scala 126:16]
  assign m_523_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_523_io_x2 = r_1469; // @[MUL.scala 104:13]
  assign m_523_io_x3 = r_1470; // @[MUL.scala 105:13]
  assign m_524_io_x1 = r_1471; // @[MUL.scala 103:13]
  assign m_524_io_x2 = r_1472; // @[MUL.scala 104:13]
  assign m_524_io_x3 = r_1473; // @[MUL.scala 105:13]
  assign m_525_io_x1 = r_1474; // @[MUL.scala 103:13]
  assign m_525_io_x2 = r_1475; // @[MUL.scala 104:13]
  assign m_525_io_x3 = r_1476; // @[MUL.scala 105:13]
  assign m_526_io_x1 = r_1477; // @[MUL.scala 103:13]
  assign m_526_io_x2 = r_1478; // @[MUL.scala 104:13]
  assign m_526_io_x3 = r_1479; // @[MUL.scala 105:13]
  assign m_527_io_x1 = r_1480; // @[MUL.scala 103:13]
  assign m_527_io_x2 = r_1481; // @[MUL.scala 104:13]
  assign m_527_io_x3 = r_1482; // @[MUL.scala 105:13]
  assign m_528_io_x1 = r_1483; // @[MUL.scala 103:13]
  assign m_528_io_x2 = r_1484; // @[MUL.scala 104:13]
  assign m_528_io_x3 = r_1485; // @[MUL.scala 105:13]
  assign m_529_io_x1 = r_1486; // @[MUL.scala 103:13]
  assign m_529_io_x2 = r_1487; // @[MUL.scala 104:13]
  assign m_529_io_x3 = r_1488; // @[MUL.scala 105:13]
  assign m_530_io_x1 = r_1489; // @[MUL.scala 103:13]
  assign m_530_io_x2 = r_1490; // @[MUL.scala 104:13]
  assign m_530_io_x3 = r_1491; // @[MUL.scala 105:13]
  assign m_531_io_x1 = r_1492; // @[MUL.scala 103:13]
  assign m_531_io_x2 = r_1493; // @[MUL.scala 104:13]
  assign m_531_io_x3 = r_1494; // @[MUL.scala 105:13]
  assign m_532_io_in_0 = r_1495; // @[MUL.scala 125:16]
  assign m_532_io_in_1 = r_1496; // @[MUL.scala 126:16]
  assign m_533_io_x1 = r_1497; // @[MUL.scala 103:13]
  assign m_533_io_x2 = r_1498; // @[MUL.scala 104:13]
  assign m_533_io_x3 = r_1499; // @[MUL.scala 105:13]
  assign m_534_io_x1 = r_1500; // @[MUL.scala 103:13]
  assign m_534_io_x2 = r_1501; // @[MUL.scala 104:13]
  assign m_534_io_x3 = r_1502; // @[MUL.scala 105:13]
  assign m_535_io_x1 = r_1503; // @[MUL.scala 103:13]
  assign m_535_io_x2 = r_1504; // @[MUL.scala 104:13]
  assign m_535_io_x3 = r_1505; // @[MUL.scala 105:13]
  assign m_536_io_x1 = r_1506; // @[MUL.scala 103:13]
  assign m_536_io_x2 = r_1507; // @[MUL.scala 104:13]
  assign m_536_io_x3 = r_1508; // @[MUL.scala 105:13]
  assign m_537_io_x1 = r_1509; // @[MUL.scala 103:13]
  assign m_537_io_x2 = r_1510; // @[MUL.scala 104:13]
  assign m_537_io_x3 = r_1511; // @[MUL.scala 105:13]
  assign m_538_io_x1 = r_1512; // @[MUL.scala 103:13]
  assign m_538_io_x2 = r_1513; // @[MUL.scala 104:13]
  assign m_538_io_x3 = r_1514; // @[MUL.scala 105:13]
  assign m_539_io_x1 = r_1515; // @[MUL.scala 103:13]
  assign m_539_io_x2 = r_1516; // @[MUL.scala 104:13]
  assign m_539_io_x3 = r_1517; // @[MUL.scala 105:13]
  assign m_540_io_x1 = r_1518; // @[MUL.scala 103:13]
  assign m_540_io_x2 = r_1519; // @[MUL.scala 104:13]
  assign m_540_io_x3 = r_1520; // @[MUL.scala 105:13]
  assign m_541_io_x1 = r_1521; // @[MUL.scala 103:13]
  assign m_541_io_x2 = r_1522; // @[MUL.scala 104:13]
  assign m_541_io_x3 = r_1523; // @[MUL.scala 105:13]
  assign m_542_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_542_io_x2 = r_1526; // @[MUL.scala 104:13]
  assign m_542_io_x3 = r_1527; // @[MUL.scala 105:13]
  assign m_543_io_x1 = r_1528; // @[MUL.scala 103:13]
  assign m_543_io_x2 = r_1529; // @[MUL.scala 104:13]
  assign m_543_io_x3 = r_1530; // @[MUL.scala 105:13]
  assign m_544_io_x1 = r_1531; // @[MUL.scala 103:13]
  assign m_544_io_x2 = r_1532; // @[MUL.scala 104:13]
  assign m_544_io_x3 = r_1533; // @[MUL.scala 105:13]
  assign m_545_io_x1 = r_1534; // @[MUL.scala 103:13]
  assign m_545_io_x2 = r_1535; // @[MUL.scala 104:13]
  assign m_545_io_x3 = r_1536; // @[MUL.scala 105:13]
  assign m_546_io_x1 = r_1537; // @[MUL.scala 103:13]
  assign m_546_io_x2 = r_1538; // @[MUL.scala 104:13]
  assign m_546_io_x3 = r_1539; // @[MUL.scala 105:13]
  assign m_547_io_x1 = r_1540; // @[MUL.scala 103:13]
  assign m_547_io_x2 = r_1541; // @[MUL.scala 104:13]
  assign m_547_io_x3 = r_1542; // @[MUL.scala 105:13]
  assign m_548_io_x1 = r_1543; // @[MUL.scala 103:13]
  assign m_548_io_x2 = r_1544; // @[MUL.scala 104:13]
  assign m_548_io_x3 = r_1545; // @[MUL.scala 105:13]
  assign m_549_io_x1 = r_1546; // @[MUL.scala 103:13]
  assign m_549_io_x2 = r_1547; // @[MUL.scala 104:13]
  assign m_549_io_x3 = r_1548; // @[MUL.scala 105:13]
  assign m_550_io_x1 = r_1549; // @[MUL.scala 103:13]
  assign m_550_io_x2 = r_1550; // @[MUL.scala 104:13]
  assign m_550_io_x3 = r_1551; // @[MUL.scala 105:13]
  assign m_551_io_x1 = r_1553; // @[MUL.scala 103:13]
  assign m_551_io_x2 = r_1554; // @[MUL.scala 104:13]
  assign m_551_io_x3 = r_1555; // @[MUL.scala 105:13]
  assign m_552_io_x1 = r_1556; // @[MUL.scala 103:13]
  assign m_552_io_x2 = r_1557; // @[MUL.scala 104:13]
  assign m_552_io_x3 = r_1558; // @[MUL.scala 105:13]
  assign m_553_io_x1 = r_1559; // @[MUL.scala 103:13]
  assign m_553_io_x2 = r_1560; // @[MUL.scala 104:13]
  assign m_553_io_x3 = r_1561; // @[MUL.scala 105:13]
  assign m_554_io_x1 = r_1562; // @[MUL.scala 103:13]
  assign m_554_io_x2 = r_1563; // @[MUL.scala 104:13]
  assign m_554_io_x3 = r_1564; // @[MUL.scala 105:13]
  assign m_555_io_x1 = r_1565; // @[MUL.scala 103:13]
  assign m_555_io_x2 = r_1566; // @[MUL.scala 104:13]
  assign m_555_io_x3 = r_1567; // @[MUL.scala 105:13]
  assign m_556_io_x1 = r_1568; // @[MUL.scala 103:13]
  assign m_556_io_x2 = r_1569; // @[MUL.scala 104:13]
  assign m_556_io_x3 = r_1570; // @[MUL.scala 105:13]
  assign m_557_io_x1 = r_1571; // @[MUL.scala 103:13]
  assign m_557_io_x2 = r_1572; // @[MUL.scala 104:13]
  assign m_557_io_x3 = r_1573; // @[MUL.scala 105:13]
  assign m_558_io_x1 = r_1574; // @[MUL.scala 103:13]
  assign m_558_io_x2 = r_1575; // @[MUL.scala 104:13]
  assign m_558_io_x3 = r_1576; // @[MUL.scala 105:13]
  assign m_559_io_x1 = r_1577; // @[MUL.scala 103:13]
  assign m_559_io_x2 = r_1578; // @[MUL.scala 104:13]
  assign m_559_io_x3 = r_1579; // @[MUL.scala 105:13]
  assign m_560_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_560_io_x2 = r_1581; // @[MUL.scala 104:13]
  assign m_560_io_x3 = r_1582; // @[MUL.scala 105:13]
  assign m_561_io_x1 = r_1583; // @[MUL.scala 103:13]
  assign m_561_io_x2 = r_1584; // @[MUL.scala 104:13]
  assign m_561_io_x3 = r_1585; // @[MUL.scala 105:13]
  assign m_562_io_x1 = r_1586; // @[MUL.scala 103:13]
  assign m_562_io_x2 = r_1587; // @[MUL.scala 104:13]
  assign m_562_io_x3 = r_1588; // @[MUL.scala 105:13]
  assign m_563_io_x1 = r_1589; // @[MUL.scala 103:13]
  assign m_563_io_x2 = r_1590; // @[MUL.scala 104:13]
  assign m_563_io_x3 = r_1591; // @[MUL.scala 105:13]
  assign m_564_io_x1 = r_1592; // @[MUL.scala 103:13]
  assign m_564_io_x2 = r_1593; // @[MUL.scala 104:13]
  assign m_564_io_x3 = r_1594; // @[MUL.scala 105:13]
  assign m_565_io_x1 = r_1595; // @[MUL.scala 103:13]
  assign m_565_io_x2 = r_1596; // @[MUL.scala 104:13]
  assign m_565_io_x3 = r_1597; // @[MUL.scala 105:13]
  assign m_566_io_x1 = r_1598; // @[MUL.scala 103:13]
  assign m_566_io_x2 = r_1599; // @[MUL.scala 104:13]
  assign m_566_io_x3 = r_1600; // @[MUL.scala 105:13]
  assign m_567_io_x1 = r_1601; // @[MUL.scala 103:13]
  assign m_567_io_x2 = r_1602; // @[MUL.scala 104:13]
  assign m_567_io_x3 = r_1603; // @[MUL.scala 105:13]
  assign m_568_io_x1 = r_1604; // @[MUL.scala 103:13]
  assign m_568_io_x2 = r_1605; // @[MUL.scala 104:13]
  assign m_568_io_x3 = r_1606; // @[MUL.scala 105:13]
  assign m_569_io_x1 = r_1607; // @[MUL.scala 103:13]
  assign m_569_io_x2 = r_1608; // @[MUL.scala 104:13]
  assign m_569_io_x3 = r_1609; // @[MUL.scala 105:13]
  assign m_570_io_x1 = r_1610; // @[MUL.scala 103:13]
  assign m_570_io_x2 = r_1611; // @[MUL.scala 104:13]
  assign m_570_io_x3 = r_1612; // @[MUL.scala 105:13]
  assign m_571_io_x1 = r_1613; // @[MUL.scala 103:13]
  assign m_571_io_x2 = r_1614; // @[MUL.scala 104:13]
  assign m_571_io_x3 = r_1615; // @[MUL.scala 105:13]
  assign m_572_io_x1 = r_1616; // @[MUL.scala 103:13]
  assign m_572_io_x2 = r_1617; // @[MUL.scala 104:13]
  assign m_572_io_x3 = r_1618; // @[MUL.scala 105:13]
  assign m_573_io_x1 = r_1619; // @[MUL.scala 103:13]
  assign m_573_io_x2 = r_1620; // @[MUL.scala 104:13]
  assign m_573_io_x3 = r_1621; // @[MUL.scala 105:13]
  assign m_574_io_x1 = r_1622; // @[MUL.scala 103:13]
  assign m_574_io_x2 = r_1623; // @[MUL.scala 104:13]
  assign m_574_io_x3 = r_1624; // @[MUL.scala 105:13]
  assign m_575_io_x1 = r_1625; // @[MUL.scala 103:13]
  assign m_575_io_x2 = r_1626; // @[MUL.scala 104:13]
  assign m_575_io_x3 = r_1627; // @[MUL.scala 105:13]
  assign m_576_io_x1 = r_1628; // @[MUL.scala 103:13]
  assign m_576_io_x2 = r_1629; // @[MUL.scala 104:13]
  assign m_576_io_x3 = r_1630; // @[MUL.scala 105:13]
  assign m_577_io_in_0 = r_1631; // @[MUL.scala 125:16]
  assign m_577_io_in_1 = r_1632; // @[MUL.scala 126:16]
  assign m_578_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_578_io_x2 = r_1634; // @[MUL.scala 104:13]
  assign m_578_io_x3 = r_1635; // @[MUL.scala 105:13]
  assign m_579_io_x1 = r_1636; // @[MUL.scala 103:13]
  assign m_579_io_x2 = r_1637; // @[MUL.scala 104:13]
  assign m_579_io_x3 = r_1638; // @[MUL.scala 105:13]
  assign m_580_io_x1 = r_1639; // @[MUL.scala 103:13]
  assign m_580_io_x2 = r_1640; // @[MUL.scala 104:13]
  assign m_580_io_x3 = r_1641; // @[MUL.scala 105:13]
  assign m_581_io_x1 = r_1642; // @[MUL.scala 103:13]
  assign m_581_io_x2 = r_1643; // @[MUL.scala 104:13]
  assign m_581_io_x3 = r_1644; // @[MUL.scala 105:13]
  assign m_582_io_x1 = r_1645; // @[MUL.scala 103:13]
  assign m_582_io_x2 = r_1646; // @[MUL.scala 104:13]
  assign m_582_io_x3 = r_1647; // @[MUL.scala 105:13]
  assign m_583_io_x1 = r_1648; // @[MUL.scala 103:13]
  assign m_583_io_x2 = r_1649; // @[MUL.scala 104:13]
  assign m_583_io_x3 = r_1650; // @[MUL.scala 105:13]
  assign m_584_io_x1 = r_1651; // @[MUL.scala 103:13]
  assign m_584_io_x2 = r_1652; // @[MUL.scala 104:13]
  assign m_584_io_x3 = r_1653; // @[MUL.scala 105:13]
  assign m_585_io_x1 = r_1654; // @[MUL.scala 103:13]
  assign m_585_io_x2 = r_1655; // @[MUL.scala 104:13]
  assign m_585_io_x3 = r_1656; // @[MUL.scala 105:13]
  assign m_586_io_in_0 = r_1657; // @[MUL.scala 125:16]
  assign m_586_io_in_1 = r_1658; // @[MUL.scala 126:16]
  assign m_587_io_x1 = r_1659; // @[MUL.scala 103:13]
  assign m_587_io_x2 = r_1660; // @[MUL.scala 104:13]
  assign m_587_io_x3 = r_1661; // @[MUL.scala 105:13]
  assign m_588_io_x1 = r_1662; // @[MUL.scala 103:13]
  assign m_588_io_x2 = r_1663; // @[MUL.scala 104:13]
  assign m_588_io_x3 = r_1664; // @[MUL.scala 105:13]
  assign m_589_io_x1 = r_1665; // @[MUL.scala 103:13]
  assign m_589_io_x2 = r_1666; // @[MUL.scala 104:13]
  assign m_589_io_x3 = r_1667; // @[MUL.scala 105:13]
  assign m_590_io_x1 = r_1668; // @[MUL.scala 103:13]
  assign m_590_io_x2 = r_1669; // @[MUL.scala 104:13]
  assign m_590_io_x3 = r_1670; // @[MUL.scala 105:13]
  assign m_591_io_x1 = r_1671; // @[MUL.scala 103:13]
  assign m_591_io_x2 = r_1672; // @[MUL.scala 104:13]
  assign m_591_io_x3 = r_1673; // @[MUL.scala 105:13]
  assign m_592_io_x1 = r_1674; // @[MUL.scala 103:13]
  assign m_592_io_x2 = r_1675; // @[MUL.scala 104:13]
  assign m_592_io_x3 = r_1676; // @[MUL.scala 105:13]
  assign m_593_io_x1 = r_1677; // @[MUL.scala 103:13]
  assign m_593_io_x2 = r_1678; // @[MUL.scala 104:13]
  assign m_593_io_x3 = r_1679; // @[MUL.scala 105:13]
  assign m_594_io_x1 = r_1680; // @[MUL.scala 103:13]
  assign m_594_io_x2 = r_1681; // @[MUL.scala 104:13]
  assign m_594_io_x3 = r_1682; // @[MUL.scala 105:13]
  assign m_595_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_595_io_x2 = r_1685; // @[MUL.scala 104:13]
  assign m_595_io_x3 = r_1686; // @[MUL.scala 105:13]
  assign m_596_io_x1 = r_1687; // @[MUL.scala 103:13]
  assign m_596_io_x2 = r_1688; // @[MUL.scala 104:13]
  assign m_596_io_x3 = r_1689; // @[MUL.scala 105:13]
  assign m_597_io_x1 = r_1690; // @[MUL.scala 103:13]
  assign m_597_io_x2 = r_1691; // @[MUL.scala 104:13]
  assign m_597_io_x3 = r_1692; // @[MUL.scala 105:13]
  assign m_598_io_x1 = r_1693; // @[MUL.scala 103:13]
  assign m_598_io_x2 = r_1694; // @[MUL.scala 104:13]
  assign m_598_io_x3 = r_1695; // @[MUL.scala 105:13]
  assign m_599_io_x1 = r_1696; // @[MUL.scala 103:13]
  assign m_599_io_x2 = r_1697; // @[MUL.scala 104:13]
  assign m_599_io_x3 = r_1698; // @[MUL.scala 105:13]
  assign m_600_io_x1 = r_1699; // @[MUL.scala 103:13]
  assign m_600_io_x2 = r_1700; // @[MUL.scala 104:13]
  assign m_600_io_x3 = r_1701; // @[MUL.scala 105:13]
  assign m_601_io_x1 = r_1702; // @[MUL.scala 103:13]
  assign m_601_io_x2 = r_1703; // @[MUL.scala 104:13]
  assign m_601_io_x3 = r_1704; // @[MUL.scala 105:13]
  assign m_602_io_x1 = r_1705; // @[MUL.scala 103:13]
  assign m_602_io_x2 = r_1706; // @[MUL.scala 104:13]
  assign m_602_io_x3 = r_1707; // @[MUL.scala 105:13]
  assign m_603_io_x1 = r_1709; // @[MUL.scala 103:13]
  assign m_603_io_x2 = r_1710; // @[MUL.scala 104:13]
  assign m_603_io_x3 = r_1711; // @[MUL.scala 105:13]
  assign m_604_io_x1 = r_1712; // @[MUL.scala 103:13]
  assign m_604_io_x2 = r_1713; // @[MUL.scala 104:13]
  assign m_604_io_x3 = r_1714; // @[MUL.scala 105:13]
  assign m_605_io_x1 = r_1715; // @[MUL.scala 103:13]
  assign m_605_io_x2 = r_1716; // @[MUL.scala 104:13]
  assign m_605_io_x3 = r_1717; // @[MUL.scala 105:13]
  assign m_606_io_x1 = r_1718; // @[MUL.scala 103:13]
  assign m_606_io_x2 = r_1719; // @[MUL.scala 104:13]
  assign m_606_io_x3 = r_1720; // @[MUL.scala 105:13]
  assign m_607_io_x1 = r_1721; // @[MUL.scala 103:13]
  assign m_607_io_x2 = r_1722; // @[MUL.scala 104:13]
  assign m_607_io_x3 = r_1723; // @[MUL.scala 105:13]
  assign m_608_io_x1 = r_1724; // @[MUL.scala 103:13]
  assign m_608_io_x2 = r_1725; // @[MUL.scala 104:13]
  assign m_608_io_x3 = r_1726; // @[MUL.scala 105:13]
  assign m_609_io_x1 = r_1727; // @[MUL.scala 103:13]
  assign m_609_io_x2 = r_1728; // @[MUL.scala 104:13]
  assign m_609_io_x3 = r_1729; // @[MUL.scala 105:13]
  assign m_610_io_x1 = r_1730; // @[MUL.scala 103:13]
  assign m_610_io_x2 = r_1731; // @[MUL.scala 104:13]
  assign m_610_io_x3 = r_1732; // @[MUL.scala 105:13]
  assign m_611_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_611_io_x2 = r_1734; // @[MUL.scala 104:13]
  assign m_611_io_x3 = r_1735; // @[MUL.scala 105:13]
  assign m_612_io_x1 = r_1736; // @[MUL.scala 103:13]
  assign m_612_io_x2 = r_1737; // @[MUL.scala 104:13]
  assign m_612_io_x3 = r_1738; // @[MUL.scala 105:13]
  assign m_613_io_x1 = r_1739; // @[MUL.scala 103:13]
  assign m_613_io_x2 = r_1740; // @[MUL.scala 104:13]
  assign m_613_io_x3 = r_1741; // @[MUL.scala 105:13]
  assign m_614_io_x1 = r_1742; // @[MUL.scala 103:13]
  assign m_614_io_x2 = r_1743; // @[MUL.scala 104:13]
  assign m_614_io_x3 = r_1744; // @[MUL.scala 105:13]
  assign m_615_io_x1 = r_1745; // @[MUL.scala 103:13]
  assign m_615_io_x2 = r_1746; // @[MUL.scala 104:13]
  assign m_615_io_x3 = r_1747; // @[MUL.scala 105:13]
  assign m_616_io_x1 = r_1748; // @[MUL.scala 103:13]
  assign m_616_io_x2 = r_1749; // @[MUL.scala 104:13]
  assign m_616_io_x3 = r_1750; // @[MUL.scala 105:13]
  assign m_617_io_x1 = r_1751; // @[MUL.scala 103:13]
  assign m_617_io_x2 = r_1752; // @[MUL.scala 104:13]
  assign m_617_io_x3 = r_1753; // @[MUL.scala 105:13]
  assign m_618_io_x1 = r_1754; // @[MUL.scala 103:13]
  assign m_618_io_x2 = r_1755; // @[MUL.scala 104:13]
  assign m_618_io_x3 = r_1756; // @[MUL.scala 105:13]
  assign m_619_io_x1 = r_1757; // @[MUL.scala 103:13]
  assign m_619_io_x2 = r_1758; // @[MUL.scala 104:13]
  assign m_619_io_x3 = r_1759; // @[MUL.scala 105:13]
  assign m_620_io_x1 = r_1760; // @[MUL.scala 103:13]
  assign m_620_io_x2 = r_1761; // @[MUL.scala 104:13]
  assign m_620_io_x3 = r_1762; // @[MUL.scala 105:13]
  assign m_621_io_x1 = r_1763; // @[MUL.scala 103:13]
  assign m_621_io_x2 = r_1764; // @[MUL.scala 104:13]
  assign m_621_io_x3 = r_1765; // @[MUL.scala 105:13]
  assign m_622_io_x1 = r_1766; // @[MUL.scala 103:13]
  assign m_622_io_x2 = r_1767; // @[MUL.scala 104:13]
  assign m_622_io_x3 = r_1768; // @[MUL.scala 105:13]
  assign m_623_io_x1 = r_1769; // @[MUL.scala 103:13]
  assign m_623_io_x2 = r_1770; // @[MUL.scala 104:13]
  assign m_623_io_x3 = r_1771; // @[MUL.scala 105:13]
  assign m_624_io_x1 = r_1772; // @[MUL.scala 103:13]
  assign m_624_io_x2 = r_1773; // @[MUL.scala 104:13]
  assign m_624_io_x3 = r_1774; // @[MUL.scala 105:13]
  assign m_625_io_x1 = r_1775; // @[MUL.scala 103:13]
  assign m_625_io_x2 = r_1776; // @[MUL.scala 104:13]
  assign m_625_io_x3 = r_1777; // @[MUL.scala 105:13]
  assign m_626_io_in_0 = r_1778; // @[MUL.scala 125:16]
  assign m_626_io_in_1 = r_1779; // @[MUL.scala 126:16]
  assign m_627_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_627_io_x2 = r_1781; // @[MUL.scala 104:13]
  assign m_627_io_x3 = r_1782; // @[MUL.scala 105:13]
  assign m_628_io_x1 = r_1783; // @[MUL.scala 103:13]
  assign m_628_io_x2 = r_1784; // @[MUL.scala 104:13]
  assign m_628_io_x3 = r_1785; // @[MUL.scala 105:13]
  assign m_629_io_x1 = r_1786; // @[MUL.scala 103:13]
  assign m_629_io_x2 = r_1787; // @[MUL.scala 104:13]
  assign m_629_io_x3 = r_1788; // @[MUL.scala 105:13]
  assign m_630_io_x1 = r_1789; // @[MUL.scala 103:13]
  assign m_630_io_x2 = r_1790; // @[MUL.scala 104:13]
  assign m_630_io_x3 = r_1791; // @[MUL.scala 105:13]
  assign m_631_io_x1 = r_1792; // @[MUL.scala 103:13]
  assign m_631_io_x2 = r_1793; // @[MUL.scala 104:13]
  assign m_631_io_x3 = r_1794; // @[MUL.scala 105:13]
  assign m_632_io_x1 = r_1795; // @[MUL.scala 103:13]
  assign m_632_io_x2 = r_1796; // @[MUL.scala 104:13]
  assign m_632_io_x3 = r_1797; // @[MUL.scala 105:13]
  assign m_633_io_x1 = r_1798; // @[MUL.scala 103:13]
  assign m_633_io_x2 = r_1799; // @[MUL.scala 104:13]
  assign m_633_io_x3 = r_1800; // @[MUL.scala 105:13]
  assign m_634_io_in_0 = r_1801; // @[MUL.scala 125:16]
  assign m_634_io_in_1 = r_1802; // @[MUL.scala 126:16]
  assign m_635_io_x1 = r_1803; // @[MUL.scala 103:13]
  assign m_635_io_x2 = r_1804; // @[MUL.scala 104:13]
  assign m_635_io_x3 = r_1805; // @[MUL.scala 105:13]
  assign m_636_io_x1 = r_1806; // @[MUL.scala 103:13]
  assign m_636_io_x2 = r_1807; // @[MUL.scala 104:13]
  assign m_636_io_x3 = r_1808; // @[MUL.scala 105:13]
  assign m_637_io_x1 = r_1809; // @[MUL.scala 103:13]
  assign m_637_io_x2 = r_1810; // @[MUL.scala 104:13]
  assign m_637_io_x3 = r_1811; // @[MUL.scala 105:13]
  assign m_638_io_x1 = r_1812; // @[MUL.scala 103:13]
  assign m_638_io_x2 = r_1813; // @[MUL.scala 104:13]
  assign m_638_io_x3 = r_1814; // @[MUL.scala 105:13]
  assign m_639_io_x1 = r_1815; // @[MUL.scala 103:13]
  assign m_639_io_x2 = r_1816; // @[MUL.scala 104:13]
  assign m_639_io_x3 = r_1817; // @[MUL.scala 105:13]
  assign m_640_io_x1 = r_1818; // @[MUL.scala 103:13]
  assign m_640_io_x2 = r_1819; // @[MUL.scala 104:13]
  assign m_640_io_x3 = r_1820; // @[MUL.scala 105:13]
  assign m_641_io_x1 = r_1821; // @[MUL.scala 103:13]
  assign m_641_io_x2 = r_1822; // @[MUL.scala 104:13]
  assign m_641_io_x3 = r_1823; // @[MUL.scala 105:13]
  assign m_642_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_642_io_x2 = r_1826; // @[MUL.scala 104:13]
  assign m_642_io_x3 = r_1827; // @[MUL.scala 105:13]
  assign m_643_io_x1 = r_1828; // @[MUL.scala 103:13]
  assign m_643_io_x2 = r_1829; // @[MUL.scala 104:13]
  assign m_643_io_x3 = r_1830; // @[MUL.scala 105:13]
  assign m_644_io_x1 = r_1831; // @[MUL.scala 103:13]
  assign m_644_io_x2 = r_1832; // @[MUL.scala 104:13]
  assign m_644_io_x3 = r_1833; // @[MUL.scala 105:13]
  assign m_645_io_x1 = r_1834; // @[MUL.scala 103:13]
  assign m_645_io_x2 = r_1835; // @[MUL.scala 104:13]
  assign m_645_io_x3 = r_1836; // @[MUL.scala 105:13]
  assign m_646_io_x1 = r_1837; // @[MUL.scala 103:13]
  assign m_646_io_x2 = r_1838; // @[MUL.scala 104:13]
  assign m_646_io_x3 = r_1839; // @[MUL.scala 105:13]
  assign m_647_io_x1 = r_1840; // @[MUL.scala 103:13]
  assign m_647_io_x2 = r_1841; // @[MUL.scala 104:13]
  assign m_647_io_x3 = r_1842; // @[MUL.scala 105:13]
  assign m_648_io_x1 = r_1843; // @[MUL.scala 103:13]
  assign m_648_io_x2 = r_1844; // @[MUL.scala 104:13]
  assign m_648_io_x3 = r_1845; // @[MUL.scala 105:13]
  assign m_649_io_x1 = r_1847; // @[MUL.scala 103:13]
  assign m_649_io_x2 = r_1848; // @[MUL.scala 104:13]
  assign m_649_io_x3 = r_1849; // @[MUL.scala 105:13]
  assign m_650_io_x1 = r_1850; // @[MUL.scala 103:13]
  assign m_650_io_x2 = r_1851; // @[MUL.scala 104:13]
  assign m_650_io_x3 = r_1852; // @[MUL.scala 105:13]
  assign m_651_io_x1 = r_1853; // @[MUL.scala 103:13]
  assign m_651_io_x2 = r_1854; // @[MUL.scala 104:13]
  assign m_651_io_x3 = r_1855; // @[MUL.scala 105:13]
  assign m_652_io_x1 = r_1856; // @[MUL.scala 103:13]
  assign m_652_io_x2 = r_1857; // @[MUL.scala 104:13]
  assign m_652_io_x3 = r_1858; // @[MUL.scala 105:13]
  assign m_653_io_x1 = r_1859; // @[MUL.scala 103:13]
  assign m_653_io_x2 = r_1860; // @[MUL.scala 104:13]
  assign m_653_io_x3 = r_1861; // @[MUL.scala 105:13]
  assign m_654_io_x1 = r_1862; // @[MUL.scala 103:13]
  assign m_654_io_x2 = r_1863; // @[MUL.scala 104:13]
  assign m_654_io_x3 = r_1864; // @[MUL.scala 105:13]
  assign m_655_io_x1 = r_1865; // @[MUL.scala 103:13]
  assign m_655_io_x2 = r_1866; // @[MUL.scala 104:13]
  assign m_655_io_x3 = r_1867; // @[MUL.scala 105:13]
  assign m_656_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_656_io_x2 = r_1869; // @[MUL.scala 104:13]
  assign m_656_io_x3 = r_1870; // @[MUL.scala 105:13]
  assign m_657_io_x1 = r_1871; // @[MUL.scala 103:13]
  assign m_657_io_x2 = r_1872; // @[MUL.scala 104:13]
  assign m_657_io_x3 = r_1873; // @[MUL.scala 105:13]
  assign m_658_io_x1 = r_1874; // @[MUL.scala 103:13]
  assign m_658_io_x2 = r_1875; // @[MUL.scala 104:13]
  assign m_658_io_x3 = r_1876; // @[MUL.scala 105:13]
  assign m_659_io_x1 = r_1877; // @[MUL.scala 103:13]
  assign m_659_io_x2 = r_1878; // @[MUL.scala 104:13]
  assign m_659_io_x3 = r_1879; // @[MUL.scala 105:13]
  assign m_660_io_x1 = r_1880; // @[MUL.scala 103:13]
  assign m_660_io_x2 = r_1881; // @[MUL.scala 104:13]
  assign m_660_io_x3 = r_1882; // @[MUL.scala 105:13]
  assign m_661_io_x1 = r_1883; // @[MUL.scala 103:13]
  assign m_661_io_x2 = r_1884; // @[MUL.scala 104:13]
  assign m_661_io_x3 = r_1885; // @[MUL.scala 105:13]
  assign m_662_io_x1 = r_1886; // @[MUL.scala 103:13]
  assign m_662_io_x2 = r_1887; // @[MUL.scala 104:13]
  assign m_662_io_x3 = r_1888; // @[MUL.scala 105:13]
  assign m_663_io_x1 = r_1889; // @[MUL.scala 103:13]
  assign m_663_io_x2 = r_1890; // @[MUL.scala 104:13]
  assign m_663_io_x3 = r_1891; // @[MUL.scala 105:13]
  assign m_664_io_x1 = r_1892; // @[MUL.scala 103:13]
  assign m_664_io_x2 = r_1893; // @[MUL.scala 104:13]
  assign m_664_io_x3 = r_1894; // @[MUL.scala 105:13]
  assign m_665_io_x1 = r_1895; // @[MUL.scala 103:13]
  assign m_665_io_x2 = r_1896; // @[MUL.scala 104:13]
  assign m_665_io_x3 = r_1897; // @[MUL.scala 105:13]
  assign m_666_io_x1 = r_1898; // @[MUL.scala 103:13]
  assign m_666_io_x2 = r_1899; // @[MUL.scala 104:13]
  assign m_666_io_x3 = r_1900; // @[MUL.scala 105:13]
  assign m_667_io_x1 = r_1901; // @[MUL.scala 103:13]
  assign m_667_io_x2 = r_1902; // @[MUL.scala 104:13]
  assign m_667_io_x3 = r_1903; // @[MUL.scala 105:13]
  assign m_668_io_x1 = r_1904; // @[MUL.scala 103:13]
  assign m_668_io_x2 = r_1905; // @[MUL.scala 104:13]
  assign m_668_io_x3 = r_1906; // @[MUL.scala 105:13]
  assign m_669_io_in_0 = r_1907; // @[MUL.scala 125:16]
  assign m_669_io_in_1 = r_1908; // @[MUL.scala 126:16]
  assign m_670_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_670_io_x2 = r_1910; // @[MUL.scala 104:13]
  assign m_670_io_x3 = r_1911; // @[MUL.scala 105:13]
  assign m_671_io_x1 = r_1912; // @[MUL.scala 103:13]
  assign m_671_io_x2 = r_1913; // @[MUL.scala 104:13]
  assign m_671_io_x3 = r_1914; // @[MUL.scala 105:13]
  assign m_672_io_x1 = r_1915; // @[MUL.scala 103:13]
  assign m_672_io_x2 = r_1916; // @[MUL.scala 104:13]
  assign m_672_io_x3 = r_1917; // @[MUL.scala 105:13]
  assign m_673_io_x1 = r_1918; // @[MUL.scala 103:13]
  assign m_673_io_x2 = r_1919; // @[MUL.scala 104:13]
  assign m_673_io_x3 = r_1920; // @[MUL.scala 105:13]
  assign m_674_io_x1 = r_1921; // @[MUL.scala 103:13]
  assign m_674_io_x2 = r_1922; // @[MUL.scala 104:13]
  assign m_674_io_x3 = r_1923; // @[MUL.scala 105:13]
  assign m_675_io_x1 = r_1924; // @[MUL.scala 103:13]
  assign m_675_io_x2 = r_1925; // @[MUL.scala 104:13]
  assign m_675_io_x3 = r_1926; // @[MUL.scala 105:13]
  assign m_676_io_in_0 = r_1927; // @[MUL.scala 125:16]
  assign m_676_io_in_1 = r_1928; // @[MUL.scala 126:16]
  assign m_677_io_x1 = r_1929; // @[MUL.scala 103:13]
  assign m_677_io_x2 = r_1930; // @[MUL.scala 104:13]
  assign m_677_io_x3 = r_1931; // @[MUL.scala 105:13]
  assign m_678_io_x1 = r_1932; // @[MUL.scala 103:13]
  assign m_678_io_x2 = r_1933; // @[MUL.scala 104:13]
  assign m_678_io_x3 = r_1934; // @[MUL.scala 105:13]
  assign m_679_io_x1 = r_1935; // @[MUL.scala 103:13]
  assign m_679_io_x2 = r_1936; // @[MUL.scala 104:13]
  assign m_679_io_x3 = r_1937; // @[MUL.scala 105:13]
  assign m_680_io_x1 = r_1938; // @[MUL.scala 103:13]
  assign m_680_io_x2 = r_1939; // @[MUL.scala 104:13]
  assign m_680_io_x3 = r_1940; // @[MUL.scala 105:13]
  assign m_681_io_x1 = r_1941; // @[MUL.scala 103:13]
  assign m_681_io_x2 = r_1942; // @[MUL.scala 104:13]
  assign m_681_io_x3 = r_1943; // @[MUL.scala 105:13]
  assign m_682_io_x1 = r_1944; // @[MUL.scala 103:13]
  assign m_682_io_x2 = r_1945; // @[MUL.scala 104:13]
  assign m_682_io_x3 = r_1946; // @[MUL.scala 105:13]
  assign m_683_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_683_io_x2 = r_1949; // @[MUL.scala 104:13]
  assign m_683_io_x3 = r_1950; // @[MUL.scala 105:13]
  assign m_684_io_x1 = r_1951; // @[MUL.scala 103:13]
  assign m_684_io_x2 = r_1952; // @[MUL.scala 104:13]
  assign m_684_io_x3 = r_1953; // @[MUL.scala 105:13]
  assign m_685_io_x1 = r_1954; // @[MUL.scala 103:13]
  assign m_685_io_x2 = r_1955; // @[MUL.scala 104:13]
  assign m_685_io_x3 = r_1956; // @[MUL.scala 105:13]
  assign m_686_io_x1 = r_1957; // @[MUL.scala 103:13]
  assign m_686_io_x2 = r_1958; // @[MUL.scala 104:13]
  assign m_686_io_x3 = r_1959; // @[MUL.scala 105:13]
  assign m_687_io_x1 = r_1960; // @[MUL.scala 103:13]
  assign m_687_io_x2 = r_1961; // @[MUL.scala 104:13]
  assign m_687_io_x3 = r_1962; // @[MUL.scala 105:13]
  assign m_688_io_x1 = r_1963; // @[MUL.scala 103:13]
  assign m_688_io_x2 = r_1964; // @[MUL.scala 104:13]
  assign m_688_io_x3 = r_1965; // @[MUL.scala 105:13]
  assign m_689_io_x1 = r_1967; // @[MUL.scala 103:13]
  assign m_689_io_x2 = r_1968; // @[MUL.scala 104:13]
  assign m_689_io_x3 = r_1969; // @[MUL.scala 105:13]
  assign m_690_io_x1 = r_1970; // @[MUL.scala 103:13]
  assign m_690_io_x2 = r_1971; // @[MUL.scala 104:13]
  assign m_690_io_x3 = r_1972; // @[MUL.scala 105:13]
  assign m_691_io_x1 = r_1973; // @[MUL.scala 103:13]
  assign m_691_io_x2 = r_1974; // @[MUL.scala 104:13]
  assign m_691_io_x3 = r_1975; // @[MUL.scala 105:13]
  assign m_692_io_x1 = r_1976; // @[MUL.scala 103:13]
  assign m_692_io_x2 = r_1977; // @[MUL.scala 104:13]
  assign m_692_io_x3 = r_1978; // @[MUL.scala 105:13]
  assign m_693_io_x1 = r_1979; // @[MUL.scala 103:13]
  assign m_693_io_x2 = r_1980; // @[MUL.scala 104:13]
  assign m_693_io_x3 = r_1981; // @[MUL.scala 105:13]
  assign m_694_io_x1 = r_1982; // @[MUL.scala 103:13]
  assign m_694_io_x2 = r_1983; // @[MUL.scala 104:13]
  assign m_694_io_x3 = r_1984; // @[MUL.scala 105:13]
  assign m_695_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_695_io_x2 = r_1986; // @[MUL.scala 104:13]
  assign m_695_io_x3 = r_1987; // @[MUL.scala 105:13]
  assign m_696_io_x1 = r_1988; // @[MUL.scala 103:13]
  assign m_696_io_x2 = r_1989; // @[MUL.scala 104:13]
  assign m_696_io_x3 = r_1990; // @[MUL.scala 105:13]
  assign m_697_io_x1 = r_1991; // @[MUL.scala 103:13]
  assign m_697_io_x2 = r_1992; // @[MUL.scala 104:13]
  assign m_697_io_x3 = r_1993; // @[MUL.scala 105:13]
  assign m_698_io_x1 = r_1994; // @[MUL.scala 103:13]
  assign m_698_io_x2 = r_1995; // @[MUL.scala 104:13]
  assign m_698_io_x3 = r_1996; // @[MUL.scala 105:13]
  assign m_699_io_x1 = r_1997; // @[MUL.scala 103:13]
  assign m_699_io_x2 = r_1998; // @[MUL.scala 104:13]
  assign m_699_io_x3 = r_1999; // @[MUL.scala 105:13]
  assign m_700_io_x1 = r_2000; // @[MUL.scala 103:13]
  assign m_700_io_x2 = r_2001; // @[MUL.scala 104:13]
  assign m_700_io_x3 = r_2002; // @[MUL.scala 105:13]
  assign m_701_io_x1 = r_2003; // @[MUL.scala 103:13]
  assign m_701_io_x2 = r_2004; // @[MUL.scala 104:13]
  assign m_701_io_x3 = r_2005; // @[MUL.scala 105:13]
  assign m_702_io_x1 = r_2006; // @[MUL.scala 103:13]
  assign m_702_io_x2 = r_2007; // @[MUL.scala 104:13]
  assign m_702_io_x3 = r_2008; // @[MUL.scala 105:13]
  assign m_703_io_x1 = r_2009; // @[MUL.scala 103:13]
  assign m_703_io_x2 = r_2010; // @[MUL.scala 104:13]
  assign m_703_io_x3 = r_2011; // @[MUL.scala 105:13]
  assign m_704_io_x1 = r_2012; // @[MUL.scala 103:13]
  assign m_704_io_x2 = r_2013; // @[MUL.scala 104:13]
  assign m_704_io_x3 = r_2014; // @[MUL.scala 105:13]
  assign m_705_io_x1 = r_2015; // @[MUL.scala 103:13]
  assign m_705_io_x2 = r_2016; // @[MUL.scala 104:13]
  assign m_705_io_x3 = r_2017; // @[MUL.scala 105:13]
  assign m_706_io_in_0 = r_2018; // @[MUL.scala 125:16]
  assign m_706_io_in_1 = r_2019; // @[MUL.scala 126:16]
  assign m_707_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_707_io_x2 = r_2021; // @[MUL.scala 104:13]
  assign m_707_io_x3 = r_2022; // @[MUL.scala 105:13]
  assign m_708_io_x1 = r_2023; // @[MUL.scala 103:13]
  assign m_708_io_x2 = r_2024; // @[MUL.scala 104:13]
  assign m_708_io_x3 = r_2025; // @[MUL.scala 105:13]
  assign m_709_io_x1 = r_2026; // @[MUL.scala 103:13]
  assign m_709_io_x2 = r_2027; // @[MUL.scala 104:13]
  assign m_709_io_x3 = r_2028; // @[MUL.scala 105:13]
  assign m_710_io_x1 = r_2029; // @[MUL.scala 103:13]
  assign m_710_io_x2 = r_2030; // @[MUL.scala 104:13]
  assign m_710_io_x3 = r_2031; // @[MUL.scala 105:13]
  assign m_711_io_x1 = r_2032; // @[MUL.scala 103:13]
  assign m_711_io_x2 = r_2033; // @[MUL.scala 104:13]
  assign m_711_io_x3 = r_2034; // @[MUL.scala 105:13]
  assign m_712_io_in_0 = r_2035; // @[MUL.scala 125:16]
  assign m_712_io_in_1 = r_2036; // @[MUL.scala 126:16]
  assign m_713_io_x1 = r_2037; // @[MUL.scala 103:13]
  assign m_713_io_x2 = r_2038; // @[MUL.scala 104:13]
  assign m_713_io_x3 = r_2039; // @[MUL.scala 105:13]
  assign m_714_io_x1 = r_2040; // @[MUL.scala 103:13]
  assign m_714_io_x2 = r_2041; // @[MUL.scala 104:13]
  assign m_714_io_x3 = r_2042; // @[MUL.scala 105:13]
  assign m_715_io_x1 = r_2043; // @[MUL.scala 103:13]
  assign m_715_io_x2 = r_2044; // @[MUL.scala 104:13]
  assign m_715_io_x3 = r_2045; // @[MUL.scala 105:13]
  assign m_716_io_x1 = r_2046; // @[MUL.scala 103:13]
  assign m_716_io_x2 = r_2047; // @[MUL.scala 104:13]
  assign m_716_io_x3 = r_2048; // @[MUL.scala 105:13]
  assign m_717_io_x1 = r_2049; // @[MUL.scala 103:13]
  assign m_717_io_x2 = r_2050; // @[MUL.scala 104:13]
  assign m_717_io_x3 = r_2051; // @[MUL.scala 105:13]
  assign m_718_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_718_io_x2 = r_2054; // @[MUL.scala 104:13]
  assign m_718_io_x3 = r_2055; // @[MUL.scala 105:13]
  assign m_719_io_x1 = r_2056; // @[MUL.scala 103:13]
  assign m_719_io_x2 = r_2057; // @[MUL.scala 104:13]
  assign m_719_io_x3 = r_2058; // @[MUL.scala 105:13]
  assign m_720_io_x1 = r_2059; // @[MUL.scala 103:13]
  assign m_720_io_x2 = r_2060; // @[MUL.scala 104:13]
  assign m_720_io_x3 = r_2061; // @[MUL.scala 105:13]
  assign m_721_io_x1 = r_2062; // @[MUL.scala 103:13]
  assign m_721_io_x2 = r_2063; // @[MUL.scala 104:13]
  assign m_721_io_x3 = r_2064; // @[MUL.scala 105:13]
  assign m_722_io_x1 = r_2065; // @[MUL.scala 103:13]
  assign m_722_io_x2 = r_2066; // @[MUL.scala 104:13]
  assign m_722_io_x3 = r_2067; // @[MUL.scala 105:13]
  assign m_723_io_x1 = r_2069; // @[MUL.scala 103:13]
  assign m_723_io_x2 = r_2070; // @[MUL.scala 104:13]
  assign m_723_io_x3 = r_2071; // @[MUL.scala 105:13]
  assign m_724_io_x1 = r_2072; // @[MUL.scala 103:13]
  assign m_724_io_x2 = r_2073; // @[MUL.scala 104:13]
  assign m_724_io_x3 = r_2074; // @[MUL.scala 105:13]
  assign m_725_io_x1 = r_2075; // @[MUL.scala 103:13]
  assign m_725_io_x2 = r_2076; // @[MUL.scala 104:13]
  assign m_725_io_x3 = r_2077; // @[MUL.scala 105:13]
  assign m_726_io_x1 = r_2078; // @[MUL.scala 103:13]
  assign m_726_io_x2 = r_2079; // @[MUL.scala 104:13]
  assign m_726_io_x3 = r_2080; // @[MUL.scala 105:13]
  assign m_727_io_x1 = r_2081; // @[MUL.scala 103:13]
  assign m_727_io_x2 = r_2082; // @[MUL.scala 104:13]
  assign m_727_io_x3 = r_2083; // @[MUL.scala 105:13]
  assign m_728_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_728_io_x2 = r_2085; // @[MUL.scala 104:13]
  assign m_728_io_x3 = r_2086; // @[MUL.scala 105:13]
  assign m_729_io_x1 = r_2087; // @[MUL.scala 103:13]
  assign m_729_io_x2 = r_2088; // @[MUL.scala 104:13]
  assign m_729_io_x3 = r_2089; // @[MUL.scala 105:13]
  assign m_730_io_x1 = r_2090; // @[MUL.scala 103:13]
  assign m_730_io_x2 = r_2091; // @[MUL.scala 104:13]
  assign m_730_io_x3 = r_2092; // @[MUL.scala 105:13]
  assign m_731_io_x1 = r_2093; // @[MUL.scala 103:13]
  assign m_731_io_x2 = r_2094; // @[MUL.scala 104:13]
  assign m_731_io_x3 = r_2095; // @[MUL.scala 105:13]
  assign m_732_io_x1 = r_2096; // @[MUL.scala 103:13]
  assign m_732_io_x2 = r_2097; // @[MUL.scala 104:13]
  assign m_732_io_x3 = r_2098; // @[MUL.scala 105:13]
  assign m_733_io_x1 = r_2099; // @[MUL.scala 103:13]
  assign m_733_io_x2 = r_2100; // @[MUL.scala 104:13]
  assign m_733_io_x3 = r_2101; // @[MUL.scala 105:13]
  assign m_734_io_x1 = r_2102; // @[MUL.scala 103:13]
  assign m_734_io_x2 = r_2103; // @[MUL.scala 104:13]
  assign m_734_io_x3 = r_2104; // @[MUL.scala 105:13]
  assign m_735_io_x1 = r_2105; // @[MUL.scala 103:13]
  assign m_735_io_x2 = r_2106; // @[MUL.scala 104:13]
  assign m_735_io_x3 = r_2107; // @[MUL.scala 105:13]
  assign m_736_io_x1 = r_2108; // @[MUL.scala 103:13]
  assign m_736_io_x2 = r_2109; // @[MUL.scala 104:13]
  assign m_736_io_x3 = r_2110; // @[MUL.scala 105:13]
  assign m_737_io_in_0 = r_2111; // @[MUL.scala 125:16]
  assign m_737_io_in_1 = r_2112; // @[MUL.scala 126:16]
  assign m_738_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_738_io_x2 = r_2114; // @[MUL.scala 104:13]
  assign m_738_io_x3 = r_2115; // @[MUL.scala 105:13]
  assign m_739_io_x1 = r_2116; // @[MUL.scala 103:13]
  assign m_739_io_x2 = r_2117; // @[MUL.scala 104:13]
  assign m_739_io_x3 = r_2118; // @[MUL.scala 105:13]
  assign m_740_io_x1 = r_2119; // @[MUL.scala 103:13]
  assign m_740_io_x2 = r_2120; // @[MUL.scala 104:13]
  assign m_740_io_x3 = r_2121; // @[MUL.scala 105:13]
  assign m_741_io_x1 = r_2122; // @[MUL.scala 103:13]
  assign m_741_io_x2 = r_2123; // @[MUL.scala 104:13]
  assign m_741_io_x3 = r_2124; // @[MUL.scala 105:13]
  assign m_742_io_in_0 = r_2125; // @[MUL.scala 125:16]
  assign m_742_io_in_1 = r_2126; // @[MUL.scala 126:16]
  assign m_743_io_x1 = r_2127; // @[MUL.scala 103:13]
  assign m_743_io_x2 = r_2128; // @[MUL.scala 104:13]
  assign m_743_io_x3 = r_2129; // @[MUL.scala 105:13]
  assign m_744_io_x1 = r_2130; // @[MUL.scala 103:13]
  assign m_744_io_x2 = r_2131; // @[MUL.scala 104:13]
  assign m_744_io_x3 = r_2132; // @[MUL.scala 105:13]
  assign m_745_io_x1 = r_2133; // @[MUL.scala 103:13]
  assign m_745_io_x2 = r_2134; // @[MUL.scala 104:13]
  assign m_745_io_x3 = r_2135; // @[MUL.scala 105:13]
  assign m_746_io_x1 = r_2136; // @[MUL.scala 103:13]
  assign m_746_io_x2 = r_2137; // @[MUL.scala 104:13]
  assign m_746_io_x3 = r_2138; // @[MUL.scala 105:13]
  assign m_747_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_747_io_x2 = r_2141; // @[MUL.scala 104:13]
  assign m_747_io_x3 = r_2142; // @[MUL.scala 105:13]
  assign m_748_io_x1 = r_2143; // @[MUL.scala 103:13]
  assign m_748_io_x2 = r_2144; // @[MUL.scala 104:13]
  assign m_748_io_x3 = r_2145; // @[MUL.scala 105:13]
  assign m_749_io_x1 = r_2146; // @[MUL.scala 103:13]
  assign m_749_io_x2 = r_2147; // @[MUL.scala 104:13]
  assign m_749_io_x3 = r_2148; // @[MUL.scala 105:13]
  assign m_750_io_x1 = r_2149; // @[MUL.scala 103:13]
  assign m_750_io_x2 = r_2150; // @[MUL.scala 104:13]
  assign m_750_io_x3 = r_2151; // @[MUL.scala 105:13]
  assign m_751_io_x1 = r_2153; // @[MUL.scala 103:13]
  assign m_751_io_x2 = r_2154; // @[MUL.scala 104:13]
  assign m_751_io_x3 = r_2155; // @[MUL.scala 105:13]
  assign m_752_io_x1 = r_2156; // @[MUL.scala 103:13]
  assign m_752_io_x2 = r_2157; // @[MUL.scala 104:13]
  assign m_752_io_x3 = r_2158; // @[MUL.scala 105:13]
  assign m_753_io_x1 = r_2159; // @[MUL.scala 103:13]
  assign m_753_io_x2 = r_2160; // @[MUL.scala 104:13]
  assign m_753_io_x3 = r_2161; // @[MUL.scala 105:13]
  assign m_754_io_x1 = r_2162; // @[MUL.scala 103:13]
  assign m_754_io_x2 = r_2163; // @[MUL.scala 104:13]
  assign m_754_io_x3 = r_2164; // @[MUL.scala 105:13]
  assign m_755_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_755_io_x2 = r_2166; // @[MUL.scala 104:13]
  assign m_755_io_x3 = r_2167; // @[MUL.scala 105:13]
  assign m_756_io_x1 = r_2168; // @[MUL.scala 103:13]
  assign m_756_io_x2 = r_2169; // @[MUL.scala 104:13]
  assign m_756_io_x3 = r_2170; // @[MUL.scala 105:13]
  assign m_757_io_x1 = r_2171; // @[MUL.scala 103:13]
  assign m_757_io_x2 = r_2172; // @[MUL.scala 104:13]
  assign m_757_io_x3 = r_2173; // @[MUL.scala 105:13]
  assign m_758_io_x1 = r_2174; // @[MUL.scala 103:13]
  assign m_758_io_x2 = r_2175; // @[MUL.scala 104:13]
  assign m_758_io_x3 = r_2176; // @[MUL.scala 105:13]
  assign m_759_io_x1 = r_2177; // @[MUL.scala 103:13]
  assign m_759_io_x2 = r_2178; // @[MUL.scala 104:13]
  assign m_759_io_x3 = r_2179; // @[MUL.scala 105:13]
  assign m_760_io_x1 = r_2180; // @[MUL.scala 103:13]
  assign m_760_io_x2 = r_2181; // @[MUL.scala 104:13]
  assign m_760_io_x3 = r_2182; // @[MUL.scala 105:13]
  assign m_761_io_x1 = r_2183; // @[MUL.scala 103:13]
  assign m_761_io_x2 = r_2184; // @[MUL.scala 104:13]
  assign m_761_io_x3 = r_2185; // @[MUL.scala 105:13]
  assign m_762_io_in_0 = r_2186; // @[MUL.scala 125:16]
  assign m_762_io_in_1 = r_2187; // @[MUL.scala 126:16]
  assign m_763_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_763_io_x2 = r_2189; // @[MUL.scala 104:13]
  assign m_763_io_x3 = r_2190; // @[MUL.scala 105:13]
  assign m_764_io_x1 = r_2191; // @[MUL.scala 103:13]
  assign m_764_io_x2 = r_2192; // @[MUL.scala 104:13]
  assign m_764_io_x3 = r_2193; // @[MUL.scala 105:13]
  assign m_765_io_x1 = r_2194; // @[MUL.scala 103:13]
  assign m_765_io_x2 = r_2195; // @[MUL.scala 104:13]
  assign m_765_io_x3 = r_2196; // @[MUL.scala 105:13]
  assign m_766_io_in_0 = r_2197; // @[MUL.scala 125:16]
  assign m_766_io_in_1 = r_2198; // @[MUL.scala 126:16]
  assign m_767_io_x1 = r_2199; // @[MUL.scala 103:13]
  assign m_767_io_x2 = r_2200; // @[MUL.scala 104:13]
  assign m_767_io_x3 = r_2201; // @[MUL.scala 105:13]
  assign m_768_io_x1 = r_2202; // @[MUL.scala 103:13]
  assign m_768_io_x2 = r_2203; // @[MUL.scala 104:13]
  assign m_768_io_x3 = r_2204; // @[MUL.scala 105:13]
  assign m_769_io_x1 = r_2205; // @[MUL.scala 103:13]
  assign m_769_io_x2 = r_2206; // @[MUL.scala 104:13]
  assign m_769_io_x3 = r_2207; // @[MUL.scala 105:13]
  assign m_770_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_770_io_x2 = r_2210; // @[MUL.scala 104:13]
  assign m_770_io_x3 = r_2211; // @[MUL.scala 105:13]
  assign m_771_io_x1 = r_2212; // @[MUL.scala 103:13]
  assign m_771_io_x2 = r_2213; // @[MUL.scala 104:13]
  assign m_771_io_x3 = r_2214; // @[MUL.scala 105:13]
  assign m_772_io_x1 = r_2215; // @[MUL.scala 103:13]
  assign m_772_io_x2 = r_2216; // @[MUL.scala 104:13]
  assign m_772_io_x3 = r_2217; // @[MUL.scala 105:13]
  assign m_773_io_x1 = r_2219; // @[MUL.scala 103:13]
  assign m_773_io_x2 = r_2220; // @[MUL.scala 104:13]
  assign m_773_io_x3 = r_2221; // @[MUL.scala 105:13]
  assign m_774_io_x1 = r_2222; // @[MUL.scala 103:13]
  assign m_774_io_x2 = r_2223; // @[MUL.scala 104:13]
  assign m_774_io_x3 = r_2224; // @[MUL.scala 105:13]
  assign m_775_io_x1 = r_2225; // @[MUL.scala 103:13]
  assign m_775_io_x2 = r_2226; // @[MUL.scala 104:13]
  assign m_775_io_x3 = r_2227; // @[MUL.scala 105:13]
  assign m_776_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_776_io_x2 = r_2229; // @[MUL.scala 104:13]
  assign m_776_io_x3 = r_2230; // @[MUL.scala 105:13]
  assign m_777_io_x1 = r_2231; // @[MUL.scala 103:13]
  assign m_777_io_x2 = r_2232; // @[MUL.scala 104:13]
  assign m_777_io_x3 = r_2233; // @[MUL.scala 105:13]
  assign m_778_io_x1 = r_2234; // @[MUL.scala 103:13]
  assign m_778_io_x2 = r_2235; // @[MUL.scala 104:13]
  assign m_778_io_x3 = r_2236; // @[MUL.scala 105:13]
  assign m_779_io_x1 = r_2237; // @[MUL.scala 103:13]
  assign m_779_io_x2 = r_2238; // @[MUL.scala 104:13]
  assign m_779_io_x3 = r_2239; // @[MUL.scala 105:13]
  assign m_780_io_x1 = r_2240; // @[MUL.scala 103:13]
  assign m_780_io_x2 = r_2241; // @[MUL.scala 104:13]
  assign m_780_io_x3 = r_2242; // @[MUL.scala 105:13]
  assign m_781_io_in_0 = r_2243; // @[MUL.scala 125:16]
  assign m_781_io_in_1 = r_2244; // @[MUL.scala 126:16]
  assign m_782_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_782_io_x2 = r_2246; // @[MUL.scala 104:13]
  assign m_782_io_x3 = r_2247; // @[MUL.scala 105:13]
  assign m_783_io_x1 = r_2248; // @[MUL.scala 103:13]
  assign m_783_io_x2 = r_2249; // @[MUL.scala 104:13]
  assign m_783_io_x3 = r_2250; // @[MUL.scala 105:13]
  assign m_784_io_in_0 = r_2251; // @[MUL.scala 125:16]
  assign m_784_io_in_1 = r_2252; // @[MUL.scala 126:16]
  assign m_785_io_x1 = r_2253; // @[MUL.scala 103:13]
  assign m_785_io_x2 = r_2254; // @[MUL.scala 104:13]
  assign m_785_io_x3 = r_2255; // @[MUL.scala 105:13]
  assign m_786_io_x1 = r_2256; // @[MUL.scala 103:13]
  assign m_786_io_x2 = r_2257; // @[MUL.scala 104:13]
  assign m_786_io_x3 = r_2258; // @[MUL.scala 105:13]
  assign m_787_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_787_io_x2 = r_2261; // @[MUL.scala 104:13]
  assign m_787_io_x3 = r_2262; // @[MUL.scala 105:13]
  assign m_788_io_x1 = r_2263; // @[MUL.scala 103:13]
  assign m_788_io_x2 = r_2264; // @[MUL.scala 104:13]
  assign m_788_io_x3 = r_2265; // @[MUL.scala 105:13]
  assign m_789_io_x1 = r_2267; // @[MUL.scala 103:13]
  assign m_789_io_x2 = r_2268; // @[MUL.scala 104:13]
  assign m_789_io_x3 = r_2269; // @[MUL.scala 105:13]
  assign m_790_io_x1 = r_2270; // @[MUL.scala 103:13]
  assign m_790_io_x2 = r_2271; // @[MUL.scala 104:13]
  assign m_790_io_x3 = r_2272; // @[MUL.scala 105:13]
  assign m_791_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_791_io_x2 = r_2274; // @[MUL.scala 104:13]
  assign m_791_io_x3 = r_2275; // @[MUL.scala 105:13]
  assign m_792_io_x1 = r_2276; // @[MUL.scala 103:13]
  assign m_792_io_x2 = r_2277; // @[MUL.scala 104:13]
  assign m_792_io_x3 = r_2278; // @[MUL.scala 105:13]
  assign m_793_io_x1 = r_2279; // @[MUL.scala 103:13]
  assign m_793_io_x2 = r_2280; // @[MUL.scala 104:13]
  assign m_793_io_x3 = r_2281; // @[MUL.scala 105:13]
  assign m_794_io_in_0 = r_2282; // @[MUL.scala 125:16]
  assign m_794_io_in_1 = r_2283; // @[MUL.scala 126:16]
  assign m_795_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_795_io_x2 = r_2285; // @[MUL.scala 104:13]
  assign m_795_io_x3 = r_2286; // @[MUL.scala 105:13]
  assign m_796_io_in_0 = r_2287; // @[MUL.scala 125:16]
  assign m_796_io_in_1 = r_2288; // @[MUL.scala 126:16]
  assign m_797_io_x1 = r_2289; // @[MUL.scala 103:13]
  assign m_797_io_x2 = r_2290; // @[MUL.scala 104:13]
  assign m_797_io_x3 = r_2291; // @[MUL.scala 105:13]
  assign m_798_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_798_io_x2 = r_2294; // @[MUL.scala 104:13]
  assign m_798_io_x3 = r_2295; // @[MUL.scala 105:13]
  assign m_799_io_x1 = r_2297; // @[MUL.scala 103:13]
  assign m_799_io_x2 = r_2298; // @[MUL.scala 104:13]
  assign m_799_io_x3 = r_2299; // @[MUL.scala 105:13]
  assign m_800_io_x1 = 1'h1; // @[MUL.scala 103:13]
  assign m_800_io_x2 = r_2301; // @[MUL.scala 104:13]
  assign m_800_io_x3 = r_2302; // @[MUL.scala 105:13]
  assign m_801_io_in_0 = r_2303; // @[MUL.scala 125:16]
  assign m_801_io_in_1 = r_2304; // @[MUL.scala 126:16]
  assign m_802_io_in_0 = 1'h1; // @[MUL.scala 125:16]
  assign m_802_io_in_1 = r_2306; // @[MUL.scala 126:16]
  assign m_803_io_in_0 = m_34_io_out_0; // @[MUL.scala 125:16]
  assign m_803_io_in_1 = m_33_io_out_1; // @[MUL.scala 126:16]
  assign m_804_io_in_0 = m_35_io_s; // @[MUL.scala 252:21]
  assign m_804_io_in_1 = m_34_io_out_1; // @[MUL.scala 126:16]
  assign m_805_io_in_0 = m_36_io_s; // @[MUL.scala 252:21]
  assign m_805_io_in_1 = m_35_io_cout; // @[MUL.scala 253:22]
  assign m_806_io_x1 = m_37_io_s; // @[MUL.scala 252:21]
  assign m_806_io_x2 = m_36_io_cout; // @[MUL.scala 253:22]
  assign m_806_io_x3 = r_13; // @[MUL.scala 105:13]
  assign m_807_io_x1 = m_38_io_s; // @[MUL.scala 252:21]
  assign m_807_io_x2 = m_37_io_cout; // @[MUL.scala 253:22]
  assign m_807_io_x3 = r_17; // @[MUL.scala 105:13]
  assign m_808_io_x1 = m_39_io_s; // @[MUL.scala 252:21]
  assign m_808_io_x2 = m_38_io_cout; // @[MUL.scala 253:22]
  assign m_808_io_x3 = m_40_io_out_0; // @[MUL.scala 105:13]
  assign m_809_io_x1 = m_41_io_s; // @[MUL.scala 252:21]
  assign m_809_io_x2 = m_39_io_cout; // @[MUL.scala 253:22]
  assign m_809_io_x3 = m_42_io_out_0; // @[MUL.scala 105:13]
  assign m_810_io_x1 = m_43_io_s; // @[MUL.scala 252:21]
  assign m_810_io_x2 = m_41_io_cout; // @[MUL.scala 253:22]
  assign m_810_io_x3 = m_44_io_s; // @[MUL.scala 252:21]
  assign m_811_io_x1 = m_45_io_s; // @[MUL.scala 252:21]
  assign m_811_io_x2 = m_43_io_cout; // @[MUL.scala 253:22]
  assign m_811_io_x3 = m_46_io_s; // @[MUL.scala 252:21]
  assign m_812_io_x1 = m_47_io_s; // @[MUL.scala 252:21]
  assign m_812_io_x2 = m_45_io_cout; // @[MUL.scala 253:22]
  assign m_812_io_x3 = m_48_io_s; // @[MUL.scala 252:21]
  assign m_813_io_in_0 = m_46_io_cout; // @[MUL.scala 253:22]
  assign m_813_io_in_1 = r_46; // @[MUL.scala 126:16]
  assign m_814_io_x1 = m_49_io_s; // @[MUL.scala 252:21]
  assign m_814_io_x2 = m_47_io_cout; // @[MUL.scala 253:22]
  assign m_814_io_x3 = m_50_io_s; // @[MUL.scala 252:21]
  assign m_815_io_in_0 = m_48_io_cout; // @[MUL.scala 253:22]
  assign m_815_io_in_1 = r_53; // @[MUL.scala 126:16]
  assign m_816_io_x1 = m_51_io_s; // @[MUL.scala 252:21]
  assign m_816_io_x2 = m_49_io_cout; // @[MUL.scala 253:22]
  assign m_816_io_x3 = m_52_io_s; // @[MUL.scala 252:21]
  assign m_817_io_in_0 = m_50_io_cout; // @[MUL.scala 253:22]
  assign m_817_io_in_1 = m_53_io_out_0; // @[MUL.scala 126:16]
  assign m_818_io_x1 = m_54_io_s; // @[MUL.scala 252:21]
  assign m_818_io_x2 = m_51_io_cout; // @[MUL.scala 253:22]
  assign m_818_io_x3 = m_55_io_s; // @[MUL.scala 252:21]
  assign m_819_io_x1 = m_52_io_cout; // @[MUL.scala 253:22]
  assign m_819_io_x2 = m_56_io_out_0; // @[MUL.scala 104:13]
  assign m_819_io_x3 = m_53_io_out_1; // @[MUL.scala 105:13]
  assign m_820_io_x1 = m_57_io_s; // @[MUL.scala 252:21]
  assign m_820_io_x2 = m_54_io_cout; // @[MUL.scala 253:22]
  assign m_820_io_x3 = m_58_io_s; // @[MUL.scala 252:21]
  assign m_821_io_x1 = m_55_io_cout; // @[MUL.scala 253:22]
  assign m_821_io_x2 = m_59_io_s; // @[MUL.scala 252:21]
  assign m_821_io_x3 = m_56_io_out_1; // @[MUL.scala 105:13]
  assign m_822_io_x1 = m_60_io_s; // @[MUL.scala 252:21]
  assign m_822_io_x2 = m_57_io_cout; // @[MUL.scala 253:22]
  assign m_822_io_x3 = m_61_io_s; // @[MUL.scala 252:21]
  assign m_823_io_x1 = m_58_io_cout; // @[MUL.scala 253:22]
  assign m_823_io_x2 = m_62_io_s; // @[MUL.scala 252:21]
  assign m_823_io_x3 = m_59_io_cout; // @[MUL.scala 253:22]
  assign m_824_io_x1 = m_63_io_s; // @[MUL.scala 252:21]
  assign m_824_io_x2 = m_60_io_cout; // @[MUL.scala 253:22]
  assign m_824_io_x3 = m_64_io_s; // @[MUL.scala 252:21]
  assign m_825_io_x1 = m_61_io_cout; // @[MUL.scala 253:22]
  assign m_825_io_x2 = m_65_io_s; // @[MUL.scala 252:21]
  assign m_825_io_x3 = m_62_io_cout; // @[MUL.scala 253:22]
  assign m_826_io_x1 = m_66_io_s; // @[MUL.scala 252:21]
  assign m_826_io_x2 = m_63_io_cout; // @[MUL.scala 253:22]
  assign m_826_io_x3 = m_67_io_s; // @[MUL.scala 252:21]
  assign m_827_io_x1 = m_64_io_cout; // @[MUL.scala 253:22]
  assign m_827_io_x2 = m_68_io_s; // @[MUL.scala 252:21]
  assign m_827_io_x3 = m_65_io_cout; // @[MUL.scala 253:22]
  assign m_828_io_x1 = m_69_io_s; // @[MUL.scala 252:21]
  assign m_828_io_x2 = m_66_io_cout; // @[MUL.scala 253:22]
  assign m_828_io_x3 = m_70_io_s; // @[MUL.scala 252:21]
  assign m_829_io_x1 = m_67_io_cout; // @[MUL.scala 253:22]
  assign m_829_io_x2 = m_71_io_s; // @[MUL.scala 252:21]
  assign m_829_io_x3 = m_68_io_cout; // @[MUL.scala 253:22]
  assign m_830_io_x1 = m_73_io_s; // @[MUL.scala 252:21]
  assign m_830_io_x2 = m_69_io_cout; // @[MUL.scala 253:22]
  assign m_830_io_x3 = m_74_io_s; // @[MUL.scala 252:21]
  assign m_831_io_x1 = m_70_io_cout; // @[MUL.scala 253:22]
  assign m_831_io_x2 = m_75_io_s; // @[MUL.scala 252:21]
  assign m_831_io_x3 = m_71_io_cout; // @[MUL.scala 253:22]
  assign m_832_io_in_0 = m_76_io_out_0; // @[MUL.scala 125:16]
  assign m_832_io_in_1 = m_72_io_out_1; // @[MUL.scala 126:16]
  assign m_833_io_x1 = m_77_io_s; // @[MUL.scala 252:21]
  assign m_833_io_x2 = m_73_io_cout; // @[MUL.scala 253:22]
  assign m_833_io_x3 = m_78_io_s; // @[MUL.scala 252:21]
  assign m_834_io_x1 = m_74_io_cout; // @[MUL.scala 253:22]
  assign m_834_io_x2 = m_79_io_s; // @[MUL.scala 252:21]
  assign m_834_io_x3 = m_75_io_cout; // @[MUL.scala 253:22]
  assign m_835_io_in_0 = m_80_io_s; // @[MUL.scala 252:21]
  assign m_835_io_in_1 = m_76_io_out_1; // @[MUL.scala 126:16]
  assign m_836_io_x1 = m_81_io_s; // @[MUL.scala 252:21]
  assign m_836_io_x2 = m_77_io_cout; // @[MUL.scala 253:22]
  assign m_836_io_x3 = m_82_io_s; // @[MUL.scala 252:21]
  assign m_837_io_x1 = m_78_io_cout; // @[MUL.scala 253:22]
  assign m_837_io_x2 = m_83_io_s; // @[MUL.scala 252:21]
  assign m_837_io_x3 = m_79_io_cout; // @[MUL.scala 253:22]
  assign m_838_io_in_0 = m_84_io_s; // @[MUL.scala 252:21]
  assign m_838_io_in_1 = m_80_io_cout; // @[MUL.scala 253:22]
  assign m_839_io_x1 = m_85_io_s; // @[MUL.scala 252:21]
  assign m_839_io_x2 = m_81_io_cout; // @[MUL.scala 253:22]
  assign m_839_io_x3 = m_86_io_s; // @[MUL.scala 252:21]
  assign m_840_io_x1 = m_82_io_cout; // @[MUL.scala 253:22]
  assign m_840_io_x2 = m_87_io_s; // @[MUL.scala 252:21]
  assign m_840_io_x3 = m_83_io_cout; // @[MUL.scala 253:22]
  assign m_841_io_x1 = m_88_io_s; // @[MUL.scala 252:21]
  assign m_841_io_x2 = m_84_io_cout; // @[MUL.scala 253:22]
  assign m_841_io_x3 = r_166; // @[MUL.scala 105:13]
  assign m_842_io_x1 = m_89_io_s; // @[MUL.scala 252:21]
  assign m_842_io_x2 = m_85_io_cout; // @[MUL.scala 253:22]
  assign m_842_io_x3 = m_90_io_s; // @[MUL.scala 252:21]
  assign m_843_io_x1 = m_86_io_cout; // @[MUL.scala 253:22]
  assign m_843_io_x2 = m_91_io_s; // @[MUL.scala 252:21]
  assign m_843_io_x3 = m_87_io_cout; // @[MUL.scala 253:22]
  assign m_844_io_x1 = m_92_io_s; // @[MUL.scala 252:21]
  assign m_844_io_x2 = m_88_io_cout; // @[MUL.scala 253:22]
  assign m_844_io_x3 = r_179; // @[MUL.scala 105:13]
  assign m_845_io_x1 = m_93_io_s; // @[MUL.scala 252:21]
  assign m_845_io_x2 = m_89_io_cout; // @[MUL.scala 253:22]
  assign m_845_io_x3 = m_94_io_s; // @[MUL.scala 252:21]
  assign m_846_io_x1 = m_90_io_cout; // @[MUL.scala 253:22]
  assign m_846_io_x2 = m_95_io_s; // @[MUL.scala 252:21]
  assign m_846_io_x3 = m_91_io_cout; // @[MUL.scala 253:22]
  assign m_847_io_x1 = m_96_io_s; // @[MUL.scala 252:21]
  assign m_847_io_x2 = m_92_io_cout; // @[MUL.scala 253:22]
  assign m_847_io_x3 = m_97_io_out_0; // @[MUL.scala 105:13]
  assign m_848_io_x1 = m_98_io_s; // @[MUL.scala 252:21]
  assign m_848_io_x2 = m_93_io_cout; // @[MUL.scala 253:22]
  assign m_848_io_x3 = m_99_io_s; // @[MUL.scala 252:21]
  assign m_849_io_x1 = m_94_io_cout; // @[MUL.scala 253:22]
  assign m_849_io_x2 = m_100_io_s; // @[MUL.scala 252:21]
  assign m_849_io_x3 = m_95_io_cout; // @[MUL.scala 253:22]
  assign m_850_io_x1 = m_101_io_s; // @[MUL.scala 252:21]
  assign m_850_io_x2 = m_96_io_cout; // @[MUL.scala 253:22]
  assign m_850_io_x3 = m_102_io_out_0; // @[MUL.scala 105:13]
  assign m_851_io_x1 = m_103_io_s; // @[MUL.scala 252:21]
  assign m_851_io_x2 = m_98_io_cout; // @[MUL.scala 253:22]
  assign m_851_io_x3 = m_104_io_s; // @[MUL.scala 252:21]
  assign m_852_io_x1 = m_99_io_cout; // @[MUL.scala 253:22]
  assign m_852_io_x2 = m_105_io_s; // @[MUL.scala 252:21]
  assign m_852_io_x3 = m_100_io_cout; // @[MUL.scala 253:22]
  assign m_853_io_x1 = m_106_io_s; // @[MUL.scala 252:21]
  assign m_853_io_x2 = m_101_io_cout; // @[MUL.scala 253:22]
  assign m_853_io_x3 = m_107_io_s; // @[MUL.scala 252:21]
  assign m_854_io_x1 = m_108_io_s; // @[MUL.scala 252:21]
  assign m_854_io_x2 = m_103_io_cout; // @[MUL.scala 253:22]
  assign m_854_io_x3 = m_109_io_s; // @[MUL.scala 252:21]
  assign m_855_io_x1 = m_104_io_cout; // @[MUL.scala 253:22]
  assign m_855_io_x2 = m_110_io_s; // @[MUL.scala 252:21]
  assign m_855_io_x3 = m_105_io_cout; // @[MUL.scala 253:22]
  assign m_856_io_x1 = m_111_io_s; // @[MUL.scala 252:21]
  assign m_856_io_x2 = m_106_io_cout; // @[MUL.scala 253:22]
  assign m_856_io_x3 = m_112_io_s; // @[MUL.scala 252:21]
  assign m_857_io_x1 = m_113_io_s; // @[MUL.scala 252:21]
  assign m_857_io_x2 = m_108_io_cout; // @[MUL.scala 253:22]
  assign m_857_io_x3 = m_114_io_s; // @[MUL.scala 252:21]
  assign m_858_io_x1 = m_109_io_cout; // @[MUL.scala 253:22]
  assign m_858_io_x2 = m_115_io_s; // @[MUL.scala 252:21]
  assign m_858_io_x3 = m_110_io_cout; // @[MUL.scala 253:22]
  assign m_859_io_x1 = m_116_io_s; // @[MUL.scala 252:21]
  assign m_859_io_x2 = m_111_io_cout; // @[MUL.scala 253:22]
  assign m_859_io_x3 = m_117_io_s; // @[MUL.scala 252:21]
  assign m_860_io_in_0 = m_112_io_cout; // @[MUL.scala 253:22]
  assign m_860_io_in_1 = r_253; // @[MUL.scala 126:16]
  assign m_861_io_x1 = m_118_io_s; // @[MUL.scala 252:21]
  assign m_861_io_x2 = m_113_io_cout; // @[MUL.scala 253:22]
  assign m_861_io_x3 = m_119_io_s; // @[MUL.scala 252:21]
  assign m_862_io_x1 = m_114_io_cout; // @[MUL.scala 253:22]
  assign m_862_io_x2 = m_120_io_s; // @[MUL.scala 252:21]
  assign m_862_io_x3 = m_115_io_cout; // @[MUL.scala 253:22]
  assign m_863_io_x1 = m_121_io_s; // @[MUL.scala 252:21]
  assign m_863_io_x2 = m_116_io_cout; // @[MUL.scala 253:22]
  assign m_863_io_x3 = m_122_io_s; // @[MUL.scala 252:21]
  assign m_864_io_in_0 = m_117_io_cout; // @[MUL.scala 253:22]
  assign m_864_io_in_1 = r_269; // @[MUL.scala 126:16]
  assign m_865_io_x1 = m_123_io_s; // @[MUL.scala 252:21]
  assign m_865_io_x2 = m_118_io_cout; // @[MUL.scala 253:22]
  assign m_865_io_x3 = m_124_io_s; // @[MUL.scala 252:21]
  assign m_866_io_x1 = m_119_io_cout; // @[MUL.scala 253:22]
  assign m_866_io_x2 = m_125_io_s; // @[MUL.scala 252:21]
  assign m_866_io_x3 = m_120_io_cout; // @[MUL.scala 253:22]
  assign m_867_io_x1 = m_126_io_s; // @[MUL.scala 252:21]
  assign m_867_io_x2 = m_121_io_cout; // @[MUL.scala 253:22]
  assign m_867_io_x3 = m_127_io_s; // @[MUL.scala 252:21]
  assign m_868_io_in_0 = m_122_io_cout; // @[MUL.scala 253:22]
  assign m_868_io_in_1 = m_128_io_out_0; // @[MUL.scala 126:16]
  assign m_869_io_x1 = m_129_io_s; // @[MUL.scala 252:21]
  assign m_869_io_x2 = m_123_io_cout; // @[MUL.scala 253:22]
  assign m_869_io_x3 = m_130_io_s; // @[MUL.scala 252:21]
  assign m_870_io_x1 = m_124_io_cout; // @[MUL.scala 253:22]
  assign m_870_io_x2 = m_131_io_s; // @[MUL.scala 252:21]
  assign m_870_io_x3 = m_125_io_cout; // @[MUL.scala 253:22]
  assign m_871_io_x1 = m_132_io_s; // @[MUL.scala 252:21]
  assign m_871_io_x2 = m_126_io_cout; // @[MUL.scala 253:22]
  assign m_871_io_x3 = m_133_io_s; // @[MUL.scala 252:21]
  assign m_872_io_x1 = m_127_io_cout; // @[MUL.scala 253:22]
  assign m_872_io_x2 = m_134_io_out_0; // @[MUL.scala 104:13]
  assign m_872_io_x3 = m_128_io_out_1; // @[MUL.scala 105:13]
  assign m_873_io_x1 = m_135_io_s; // @[MUL.scala 252:21]
  assign m_873_io_x2 = m_129_io_cout; // @[MUL.scala 253:22]
  assign m_873_io_x3 = m_136_io_s; // @[MUL.scala 252:21]
  assign m_874_io_x1 = m_130_io_cout; // @[MUL.scala 253:22]
  assign m_874_io_x2 = m_137_io_s; // @[MUL.scala 252:21]
  assign m_874_io_x3 = m_131_io_cout; // @[MUL.scala 253:22]
  assign m_875_io_x1 = m_138_io_s; // @[MUL.scala 252:21]
  assign m_875_io_x2 = m_132_io_cout; // @[MUL.scala 253:22]
  assign m_875_io_x3 = m_139_io_s; // @[MUL.scala 252:21]
  assign m_876_io_x1 = m_133_io_cout; // @[MUL.scala 253:22]
  assign m_876_io_x2 = m_140_io_s; // @[MUL.scala 252:21]
  assign m_876_io_x3 = m_134_io_out_1; // @[MUL.scala 105:13]
  assign m_877_io_x1 = m_141_io_s; // @[MUL.scala 252:21]
  assign m_877_io_x2 = m_135_io_cout; // @[MUL.scala 253:22]
  assign m_877_io_x3 = m_142_io_s; // @[MUL.scala 252:21]
  assign m_878_io_x1 = m_136_io_cout; // @[MUL.scala 253:22]
  assign m_878_io_x2 = m_143_io_s; // @[MUL.scala 252:21]
  assign m_878_io_x3 = m_137_io_cout; // @[MUL.scala 253:22]
  assign m_879_io_x1 = m_144_io_s; // @[MUL.scala 252:21]
  assign m_879_io_x2 = m_138_io_cout; // @[MUL.scala 253:22]
  assign m_879_io_x3 = m_145_io_s; // @[MUL.scala 252:21]
  assign m_880_io_x1 = m_139_io_cout; // @[MUL.scala 253:22]
  assign m_880_io_x2 = m_146_io_s; // @[MUL.scala 252:21]
  assign m_880_io_x3 = m_140_io_cout; // @[MUL.scala 253:22]
  assign m_881_io_x1 = m_147_io_s; // @[MUL.scala 252:21]
  assign m_881_io_x2 = m_141_io_cout; // @[MUL.scala 253:22]
  assign m_881_io_x3 = m_148_io_s; // @[MUL.scala 252:21]
  assign m_882_io_x1 = m_142_io_cout; // @[MUL.scala 253:22]
  assign m_882_io_x2 = m_149_io_s; // @[MUL.scala 252:21]
  assign m_882_io_x3 = m_143_io_cout; // @[MUL.scala 253:22]
  assign m_883_io_x1 = m_150_io_s; // @[MUL.scala 252:21]
  assign m_883_io_x2 = m_144_io_cout; // @[MUL.scala 253:22]
  assign m_883_io_x3 = m_151_io_s; // @[MUL.scala 252:21]
  assign m_884_io_x1 = m_145_io_cout; // @[MUL.scala 253:22]
  assign m_884_io_x2 = m_152_io_s; // @[MUL.scala 252:21]
  assign m_884_io_x3 = m_146_io_cout; // @[MUL.scala 253:22]
  assign m_885_io_x1 = m_153_io_s; // @[MUL.scala 252:21]
  assign m_885_io_x2 = m_147_io_cout; // @[MUL.scala 253:22]
  assign m_885_io_x3 = m_154_io_s; // @[MUL.scala 252:21]
  assign m_886_io_x1 = m_148_io_cout; // @[MUL.scala 253:22]
  assign m_886_io_x2 = m_155_io_s; // @[MUL.scala 252:21]
  assign m_886_io_x3 = m_149_io_cout; // @[MUL.scala 253:22]
  assign m_887_io_x1 = m_156_io_s; // @[MUL.scala 252:21]
  assign m_887_io_x2 = m_150_io_cout; // @[MUL.scala 253:22]
  assign m_887_io_x3 = m_157_io_s; // @[MUL.scala 252:21]
  assign m_888_io_x1 = m_151_io_cout; // @[MUL.scala 253:22]
  assign m_888_io_x2 = m_158_io_s; // @[MUL.scala 252:21]
  assign m_888_io_x3 = m_152_io_cout; // @[MUL.scala 253:22]
  assign m_889_io_x1 = m_159_io_s; // @[MUL.scala 252:21]
  assign m_889_io_x2 = m_153_io_cout; // @[MUL.scala 253:22]
  assign m_889_io_x3 = m_160_io_s; // @[MUL.scala 252:21]
  assign m_890_io_x1 = m_154_io_cout; // @[MUL.scala 253:22]
  assign m_890_io_x2 = m_161_io_s; // @[MUL.scala 252:21]
  assign m_890_io_x3 = m_155_io_cout; // @[MUL.scala 253:22]
  assign m_891_io_x1 = m_162_io_s; // @[MUL.scala 252:21]
  assign m_891_io_x2 = m_156_io_cout; // @[MUL.scala 253:22]
  assign m_891_io_x3 = m_163_io_s; // @[MUL.scala 252:21]
  assign m_892_io_x1 = m_157_io_cout; // @[MUL.scala 253:22]
  assign m_892_io_x2 = m_164_io_s; // @[MUL.scala 252:21]
  assign m_892_io_x3 = m_158_io_cout; // @[MUL.scala 253:22]
  assign m_893_io_x1 = m_166_io_s; // @[MUL.scala 252:21]
  assign m_893_io_x2 = m_159_io_cout; // @[MUL.scala 253:22]
  assign m_893_io_x3 = m_167_io_s; // @[MUL.scala 252:21]
  assign m_894_io_x1 = m_160_io_cout; // @[MUL.scala 253:22]
  assign m_894_io_x2 = m_168_io_s; // @[MUL.scala 252:21]
  assign m_894_io_x3 = m_161_io_cout; // @[MUL.scala 253:22]
  assign m_895_io_x1 = m_169_io_s; // @[MUL.scala 252:21]
  assign m_895_io_x2 = m_162_io_cout; // @[MUL.scala 253:22]
  assign m_895_io_x3 = m_170_io_s; // @[MUL.scala 252:21]
  assign m_896_io_x1 = m_163_io_cout; // @[MUL.scala 253:22]
  assign m_896_io_x2 = m_171_io_s; // @[MUL.scala 252:21]
  assign m_896_io_x3 = m_164_io_cout; // @[MUL.scala 253:22]
  assign m_897_io_in_0 = m_172_io_out_0; // @[MUL.scala 125:16]
  assign m_897_io_in_1 = m_165_io_out_1; // @[MUL.scala 126:16]
  assign m_898_io_x1 = m_173_io_s; // @[MUL.scala 252:21]
  assign m_898_io_x2 = m_166_io_cout; // @[MUL.scala 253:22]
  assign m_898_io_x3 = m_174_io_s; // @[MUL.scala 252:21]
  assign m_899_io_x1 = m_167_io_cout; // @[MUL.scala 253:22]
  assign m_899_io_x2 = m_175_io_s; // @[MUL.scala 252:21]
  assign m_899_io_x3 = m_168_io_cout; // @[MUL.scala 253:22]
  assign m_900_io_x1 = m_176_io_s; // @[MUL.scala 252:21]
  assign m_900_io_x2 = m_169_io_cout; // @[MUL.scala 253:22]
  assign m_900_io_x3 = m_177_io_s; // @[MUL.scala 252:21]
  assign m_901_io_x1 = m_170_io_cout; // @[MUL.scala 253:22]
  assign m_901_io_x2 = m_178_io_s; // @[MUL.scala 252:21]
  assign m_901_io_x3 = m_171_io_cout; // @[MUL.scala 253:22]
  assign m_902_io_in_0 = m_179_io_s; // @[MUL.scala 252:21]
  assign m_902_io_in_1 = m_172_io_out_1; // @[MUL.scala 126:16]
  assign m_903_io_x1 = m_180_io_s; // @[MUL.scala 252:21]
  assign m_903_io_x2 = m_173_io_cout; // @[MUL.scala 253:22]
  assign m_903_io_x3 = m_181_io_s; // @[MUL.scala 252:21]
  assign m_904_io_x1 = m_174_io_cout; // @[MUL.scala 253:22]
  assign m_904_io_x2 = m_182_io_s; // @[MUL.scala 252:21]
  assign m_904_io_x3 = m_175_io_cout; // @[MUL.scala 253:22]
  assign m_905_io_x1 = m_183_io_s; // @[MUL.scala 252:21]
  assign m_905_io_x2 = m_176_io_cout; // @[MUL.scala 253:22]
  assign m_905_io_x3 = m_184_io_s; // @[MUL.scala 252:21]
  assign m_906_io_x1 = m_177_io_cout; // @[MUL.scala 253:22]
  assign m_906_io_x2 = m_185_io_s; // @[MUL.scala 252:21]
  assign m_906_io_x3 = m_178_io_cout; // @[MUL.scala 253:22]
  assign m_907_io_in_0 = m_186_io_s; // @[MUL.scala 252:21]
  assign m_907_io_in_1 = m_179_io_cout; // @[MUL.scala 253:22]
  assign m_908_io_x1 = m_187_io_s; // @[MUL.scala 252:21]
  assign m_908_io_x2 = m_180_io_cout; // @[MUL.scala 253:22]
  assign m_908_io_x3 = m_188_io_s; // @[MUL.scala 252:21]
  assign m_909_io_x1 = m_181_io_cout; // @[MUL.scala 253:22]
  assign m_909_io_x2 = m_189_io_s; // @[MUL.scala 252:21]
  assign m_909_io_x3 = m_182_io_cout; // @[MUL.scala 253:22]
  assign m_910_io_x1 = m_190_io_s; // @[MUL.scala 252:21]
  assign m_910_io_x2 = m_183_io_cout; // @[MUL.scala 253:22]
  assign m_910_io_x3 = m_191_io_s; // @[MUL.scala 252:21]
  assign m_911_io_x1 = m_184_io_cout; // @[MUL.scala 253:22]
  assign m_911_io_x2 = m_192_io_s; // @[MUL.scala 252:21]
  assign m_911_io_x3 = m_185_io_cout; // @[MUL.scala 253:22]
  assign m_912_io_x1 = m_193_io_s; // @[MUL.scala 252:21]
  assign m_912_io_x2 = m_186_io_cout; // @[MUL.scala 253:22]
  assign m_912_io_x3 = r_481; // @[MUL.scala 105:13]
  assign m_913_io_x1 = m_194_io_s; // @[MUL.scala 252:21]
  assign m_913_io_x2 = m_187_io_cout; // @[MUL.scala 253:22]
  assign m_913_io_x3 = m_195_io_s; // @[MUL.scala 252:21]
  assign m_914_io_x1 = m_188_io_cout; // @[MUL.scala 253:22]
  assign m_914_io_x2 = m_196_io_s; // @[MUL.scala 252:21]
  assign m_914_io_x3 = m_189_io_cout; // @[MUL.scala 253:22]
  assign m_915_io_x1 = m_197_io_s; // @[MUL.scala 252:21]
  assign m_915_io_x2 = m_190_io_cout; // @[MUL.scala 253:22]
  assign m_915_io_x3 = m_198_io_s; // @[MUL.scala 252:21]
  assign m_916_io_x1 = m_191_io_cout; // @[MUL.scala 253:22]
  assign m_916_io_x2 = m_199_io_s; // @[MUL.scala 252:21]
  assign m_916_io_x3 = m_192_io_cout; // @[MUL.scala 253:22]
  assign m_917_io_x1 = m_200_io_s; // @[MUL.scala 252:21]
  assign m_917_io_x2 = m_193_io_cout; // @[MUL.scala 253:22]
  assign m_917_io_x3 = r_503; // @[MUL.scala 105:13]
  assign m_918_io_x1 = m_201_io_s; // @[MUL.scala 252:21]
  assign m_918_io_x2 = m_194_io_cout; // @[MUL.scala 253:22]
  assign m_918_io_x3 = m_202_io_s; // @[MUL.scala 252:21]
  assign m_919_io_x1 = m_195_io_cout; // @[MUL.scala 253:22]
  assign m_919_io_x2 = m_203_io_s; // @[MUL.scala 252:21]
  assign m_919_io_x3 = m_196_io_cout; // @[MUL.scala 253:22]
  assign m_920_io_x1 = m_204_io_s; // @[MUL.scala 252:21]
  assign m_920_io_x2 = m_197_io_cout; // @[MUL.scala 253:22]
  assign m_920_io_x3 = m_205_io_s; // @[MUL.scala 252:21]
  assign m_921_io_x1 = m_198_io_cout; // @[MUL.scala 253:22]
  assign m_921_io_x2 = m_206_io_s; // @[MUL.scala 252:21]
  assign m_921_io_x3 = m_199_io_cout; // @[MUL.scala 253:22]
  assign m_922_io_x1 = m_207_io_s; // @[MUL.scala 252:21]
  assign m_922_io_x2 = m_200_io_cout; // @[MUL.scala 253:22]
  assign m_922_io_x3 = m_208_io_out_0; // @[MUL.scala 105:13]
  assign m_923_io_x1 = m_209_io_s; // @[MUL.scala 252:21]
  assign m_923_io_x2 = m_201_io_cout; // @[MUL.scala 253:22]
  assign m_923_io_x3 = m_210_io_s; // @[MUL.scala 252:21]
  assign m_924_io_x1 = m_202_io_cout; // @[MUL.scala 253:22]
  assign m_924_io_x2 = m_211_io_s; // @[MUL.scala 252:21]
  assign m_924_io_x3 = m_203_io_cout; // @[MUL.scala 253:22]
  assign m_925_io_x1 = m_212_io_s; // @[MUL.scala 252:21]
  assign m_925_io_x2 = m_204_io_cout; // @[MUL.scala 253:22]
  assign m_925_io_x3 = m_213_io_s; // @[MUL.scala 252:21]
  assign m_926_io_x1 = m_205_io_cout; // @[MUL.scala 253:22]
  assign m_926_io_x2 = m_214_io_s; // @[MUL.scala 252:21]
  assign m_926_io_x3 = m_206_io_cout; // @[MUL.scala 253:22]
  assign m_927_io_x1 = m_215_io_s; // @[MUL.scala 252:21]
  assign m_927_io_x2 = m_207_io_cout; // @[MUL.scala 253:22]
  assign m_927_io_x3 = m_216_io_out_0; // @[MUL.scala 105:13]
  assign m_928_io_x1 = m_217_io_s; // @[MUL.scala 252:21]
  assign m_928_io_x2 = m_209_io_cout; // @[MUL.scala 253:22]
  assign m_928_io_x3 = m_218_io_s; // @[MUL.scala 252:21]
  assign m_929_io_x1 = m_210_io_cout; // @[MUL.scala 253:22]
  assign m_929_io_x2 = m_219_io_s; // @[MUL.scala 252:21]
  assign m_929_io_x3 = m_211_io_cout; // @[MUL.scala 253:22]
  assign m_930_io_x1 = m_220_io_s; // @[MUL.scala 252:21]
  assign m_930_io_x2 = m_212_io_cout; // @[MUL.scala 253:22]
  assign m_930_io_x3 = m_221_io_s; // @[MUL.scala 252:21]
  assign m_931_io_x1 = m_213_io_cout; // @[MUL.scala 253:22]
  assign m_931_io_x2 = m_222_io_s; // @[MUL.scala 252:21]
  assign m_931_io_x3 = m_214_io_cout; // @[MUL.scala 253:22]
  assign m_932_io_x1 = m_223_io_s; // @[MUL.scala 252:21]
  assign m_932_io_x2 = m_215_io_cout; // @[MUL.scala 253:22]
  assign m_932_io_x3 = m_224_io_s; // @[MUL.scala 252:21]
  assign m_933_io_x1 = m_225_io_s; // @[MUL.scala 252:21]
  assign m_933_io_x2 = m_217_io_cout; // @[MUL.scala 253:22]
  assign m_933_io_x3 = m_226_io_s; // @[MUL.scala 252:21]
  assign m_934_io_x1 = m_218_io_cout; // @[MUL.scala 253:22]
  assign m_934_io_x2 = m_227_io_s; // @[MUL.scala 252:21]
  assign m_934_io_x3 = m_219_io_cout; // @[MUL.scala 253:22]
  assign m_935_io_x1 = m_228_io_s; // @[MUL.scala 252:21]
  assign m_935_io_x2 = m_220_io_cout; // @[MUL.scala 253:22]
  assign m_935_io_x3 = m_229_io_s; // @[MUL.scala 252:21]
  assign m_936_io_x1 = m_221_io_cout; // @[MUL.scala 253:22]
  assign m_936_io_x2 = m_230_io_s; // @[MUL.scala 252:21]
  assign m_936_io_x3 = m_222_io_cout; // @[MUL.scala 253:22]
  assign m_937_io_x1 = m_231_io_s; // @[MUL.scala 252:21]
  assign m_937_io_x2 = m_223_io_cout; // @[MUL.scala 253:22]
  assign m_937_io_x3 = m_232_io_s; // @[MUL.scala 252:21]
  assign m_938_io_x1 = m_233_io_s; // @[MUL.scala 252:21]
  assign m_938_io_x2 = m_225_io_cout; // @[MUL.scala 253:22]
  assign m_938_io_x3 = m_234_io_s; // @[MUL.scala 252:21]
  assign m_939_io_x1 = m_226_io_cout; // @[MUL.scala 253:22]
  assign m_939_io_x2 = m_235_io_s; // @[MUL.scala 252:21]
  assign m_939_io_x3 = m_227_io_cout; // @[MUL.scala 253:22]
  assign m_940_io_x1 = m_236_io_s; // @[MUL.scala 252:21]
  assign m_940_io_x2 = m_228_io_cout; // @[MUL.scala 253:22]
  assign m_940_io_x3 = m_237_io_s; // @[MUL.scala 252:21]
  assign m_941_io_x1 = m_229_io_cout; // @[MUL.scala 253:22]
  assign m_941_io_x2 = m_238_io_s; // @[MUL.scala 252:21]
  assign m_941_io_x3 = m_230_io_cout; // @[MUL.scala 253:22]
  assign m_942_io_x1 = m_239_io_s; // @[MUL.scala 252:21]
  assign m_942_io_x2 = m_231_io_cout; // @[MUL.scala 253:22]
  assign m_942_io_x3 = m_240_io_s; // @[MUL.scala 252:21]
  assign m_943_io_in_0 = m_232_io_cout; // @[MUL.scala 253:22]
  assign m_943_io_in_1 = r_622; // @[MUL.scala 126:16]
  assign m_944_io_x1 = m_241_io_s; // @[MUL.scala 252:21]
  assign m_944_io_x2 = m_233_io_cout; // @[MUL.scala 253:22]
  assign m_944_io_x3 = m_242_io_s; // @[MUL.scala 252:21]
  assign m_945_io_x1 = m_234_io_cout; // @[MUL.scala 253:22]
  assign m_945_io_x2 = m_243_io_s; // @[MUL.scala 252:21]
  assign m_945_io_x3 = m_235_io_cout; // @[MUL.scala 253:22]
  assign m_946_io_x1 = m_244_io_s; // @[MUL.scala 252:21]
  assign m_946_io_x2 = m_236_io_cout; // @[MUL.scala 253:22]
  assign m_946_io_x3 = m_245_io_s; // @[MUL.scala 252:21]
  assign m_947_io_x1 = m_237_io_cout; // @[MUL.scala 253:22]
  assign m_947_io_x2 = m_246_io_s; // @[MUL.scala 252:21]
  assign m_947_io_x3 = m_238_io_cout; // @[MUL.scala 253:22]
  assign m_948_io_x1 = m_247_io_s; // @[MUL.scala 252:21]
  assign m_948_io_x2 = m_239_io_cout; // @[MUL.scala 253:22]
  assign m_948_io_x3 = m_248_io_s; // @[MUL.scala 252:21]
  assign m_949_io_in_0 = m_240_io_cout; // @[MUL.scala 253:22]
  assign m_949_io_in_1 = r_647; // @[MUL.scala 126:16]
  assign m_950_io_x1 = m_249_io_s; // @[MUL.scala 252:21]
  assign m_950_io_x2 = m_241_io_cout; // @[MUL.scala 253:22]
  assign m_950_io_x3 = m_250_io_s; // @[MUL.scala 252:21]
  assign m_951_io_x1 = m_242_io_cout; // @[MUL.scala 253:22]
  assign m_951_io_x2 = m_251_io_s; // @[MUL.scala 252:21]
  assign m_951_io_x3 = m_243_io_cout; // @[MUL.scala 253:22]
  assign m_952_io_x1 = m_252_io_s; // @[MUL.scala 252:21]
  assign m_952_io_x2 = m_244_io_cout; // @[MUL.scala 253:22]
  assign m_952_io_x3 = m_253_io_s; // @[MUL.scala 252:21]
  assign m_953_io_x1 = m_245_io_cout; // @[MUL.scala 253:22]
  assign m_953_io_x2 = m_254_io_s; // @[MUL.scala 252:21]
  assign m_953_io_x3 = m_246_io_cout; // @[MUL.scala 253:22]
  assign m_954_io_x1 = m_255_io_s; // @[MUL.scala 252:21]
  assign m_954_io_x2 = m_247_io_cout; // @[MUL.scala 253:22]
  assign m_954_io_x3 = m_256_io_s; // @[MUL.scala 252:21]
  assign m_955_io_in_0 = m_248_io_cout; // @[MUL.scala 253:22]
  assign m_955_io_in_1 = m_257_io_out_0; // @[MUL.scala 126:16]
  assign m_956_io_x1 = m_258_io_s; // @[MUL.scala 252:21]
  assign m_956_io_x2 = m_249_io_cout; // @[MUL.scala 253:22]
  assign m_956_io_x3 = m_259_io_s; // @[MUL.scala 252:21]
  assign m_957_io_x1 = m_250_io_cout; // @[MUL.scala 253:22]
  assign m_957_io_x2 = m_260_io_s; // @[MUL.scala 252:21]
  assign m_957_io_x3 = m_251_io_cout; // @[MUL.scala 253:22]
  assign m_958_io_x1 = m_261_io_s; // @[MUL.scala 252:21]
  assign m_958_io_x2 = m_252_io_cout; // @[MUL.scala 253:22]
  assign m_958_io_x3 = m_262_io_s; // @[MUL.scala 252:21]
  assign m_959_io_x1 = m_253_io_cout; // @[MUL.scala 253:22]
  assign m_959_io_x2 = m_263_io_s; // @[MUL.scala 252:21]
  assign m_959_io_x3 = m_254_io_cout; // @[MUL.scala 253:22]
  assign m_960_io_x1 = m_264_io_s; // @[MUL.scala 252:21]
  assign m_960_io_x2 = m_255_io_cout; // @[MUL.scala 253:22]
  assign m_960_io_x3 = m_265_io_s; // @[MUL.scala 252:21]
  assign m_961_io_x1 = m_256_io_cout; // @[MUL.scala 253:22]
  assign m_961_io_x2 = m_266_io_out_0; // @[MUL.scala 104:13]
  assign m_961_io_x3 = m_257_io_out_1; // @[MUL.scala 105:13]
  assign m_962_io_x1 = m_267_io_s; // @[MUL.scala 252:21]
  assign m_962_io_x2 = m_258_io_cout; // @[MUL.scala 253:22]
  assign m_962_io_x3 = m_268_io_s; // @[MUL.scala 252:21]
  assign m_963_io_x1 = m_259_io_cout; // @[MUL.scala 253:22]
  assign m_963_io_x2 = m_269_io_s; // @[MUL.scala 252:21]
  assign m_963_io_x3 = m_260_io_cout; // @[MUL.scala 253:22]
  assign m_964_io_x1 = m_270_io_s; // @[MUL.scala 252:21]
  assign m_964_io_x2 = m_261_io_cout; // @[MUL.scala 253:22]
  assign m_964_io_x3 = m_271_io_s; // @[MUL.scala 252:21]
  assign m_965_io_x1 = m_262_io_cout; // @[MUL.scala 253:22]
  assign m_965_io_x2 = m_272_io_s; // @[MUL.scala 252:21]
  assign m_965_io_x3 = m_263_io_cout; // @[MUL.scala 253:22]
  assign m_966_io_x1 = m_273_io_s; // @[MUL.scala 252:21]
  assign m_966_io_x2 = m_264_io_cout; // @[MUL.scala 253:22]
  assign m_966_io_x3 = m_274_io_s; // @[MUL.scala 252:21]
  assign m_967_io_x1 = m_265_io_cout; // @[MUL.scala 253:22]
  assign m_967_io_x2 = m_275_io_s; // @[MUL.scala 252:21]
  assign m_967_io_x3 = m_266_io_out_1; // @[MUL.scala 105:13]
  assign m_968_io_x1 = m_276_io_s; // @[MUL.scala 252:21]
  assign m_968_io_x2 = m_267_io_cout; // @[MUL.scala 253:22]
  assign m_968_io_x3 = m_277_io_s; // @[MUL.scala 252:21]
  assign m_969_io_x1 = m_268_io_cout; // @[MUL.scala 253:22]
  assign m_969_io_x2 = m_278_io_s; // @[MUL.scala 252:21]
  assign m_969_io_x3 = m_269_io_cout; // @[MUL.scala 253:22]
  assign m_970_io_x1 = m_279_io_s; // @[MUL.scala 252:21]
  assign m_970_io_x2 = m_270_io_cout; // @[MUL.scala 253:22]
  assign m_970_io_x3 = m_280_io_s; // @[MUL.scala 252:21]
  assign m_971_io_x1 = m_271_io_cout; // @[MUL.scala 253:22]
  assign m_971_io_x2 = m_281_io_s; // @[MUL.scala 252:21]
  assign m_971_io_x3 = m_272_io_cout; // @[MUL.scala 253:22]
  assign m_972_io_x1 = m_282_io_s; // @[MUL.scala 252:21]
  assign m_972_io_x2 = m_273_io_cout; // @[MUL.scala 253:22]
  assign m_972_io_x3 = m_283_io_s; // @[MUL.scala 252:21]
  assign m_973_io_x1 = m_274_io_cout; // @[MUL.scala 253:22]
  assign m_973_io_x2 = m_284_io_s; // @[MUL.scala 252:21]
  assign m_973_io_x3 = m_275_io_cout; // @[MUL.scala 253:22]
  assign m_974_io_x1 = m_285_io_s; // @[MUL.scala 252:21]
  assign m_974_io_x2 = m_276_io_cout; // @[MUL.scala 253:22]
  assign m_974_io_x3 = m_286_io_s; // @[MUL.scala 252:21]
  assign m_975_io_x1 = m_277_io_cout; // @[MUL.scala 253:22]
  assign m_975_io_x2 = m_287_io_s; // @[MUL.scala 252:21]
  assign m_975_io_x3 = m_278_io_cout; // @[MUL.scala 253:22]
  assign m_976_io_x1 = m_288_io_s; // @[MUL.scala 252:21]
  assign m_976_io_x2 = m_279_io_cout; // @[MUL.scala 253:22]
  assign m_976_io_x3 = m_289_io_s; // @[MUL.scala 252:21]
  assign m_977_io_x1 = m_280_io_cout; // @[MUL.scala 253:22]
  assign m_977_io_x2 = m_290_io_s; // @[MUL.scala 252:21]
  assign m_977_io_x3 = m_281_io_cout; // @[MUL.scala 253:22]
  assign m_978_io_x1 = m_291_io_s; // @[MUL.scala 252:21]
  assign m_978_io_x2 = m_282_io_cout; // @[MUL.scala 253:22]
  assign m_978_io_x3 = m_292_io_s; // @[MUL.scala 252:21]
  assign m_979_io_x1 = m_283_io_cout; // @[MUL.scala 253:22]
  assign m_979_io_x2 = m_293_io_s; // @[MUL.scala 252:21]
  assign m_979_io_x3 = m_284_io_cout; // @[MUL.scala 253:22]
  assign m_980_io_x1 = m_294_io_s; // @[MUL.scala 252:21]
  assign m_980_io_x2 = m_285_io_cout; // @[MUL.scala 253:22]
  assign m_980_io_x3 = m_295_io_s; // @[MUL.scala 252:21]
  assign m_981_io_x1 = m_286_io_cout; // @[MUL.scala 253:22]
  assign m_981_io_x2 = m_296_io_s; // @[MUL.scala 252:21]
  assign m_981_io_x3 = m_287_io_cout; // @[MUL.scala 253:22]
  assign m_982_io_x1 = m_297_io_s; // @[MUL.scala 252:21]
  assign m_982_io_x2 = m_288_io_cout; // @[MUL.scala 253:22]
  assign m_982_io_x3 = m_298_io_s; // @[MUL.scala 252:21]
  assign m_983_io_x1 = m_289_io_cout; // @[MUL.scala 253:22]
  assign m_983_io_x2 = m_299_io_s; // @[MUL.scala 252:21]
  assign m_983_io_x3 = m_290_io_cout; // @[MUL.scala 253:22]
  assign m_984_io_x1 = m_300_io_s; // @[MUL.scala 252:21]
  assign m_984_io_x2 = m_291_io_cout; // @[MUL.scala 253:22]
  assign m_984_io_x3 = m_301_io_s; // @[MUL.scala 252:21]
  assign m_985_io_x1 = m_292_io_cout; // @[MUL.scala 253:22]
  assign m_985_io_x2 = m_302_io_s; // @[MUL.scala 252:21]
  assign m_985_io_x3 = m_293_io_cout; // @[MUL.scala 253:22]
  assign m_986_io_x1 = m_303_io_s; // @[MUL.scala 252:21]
  assign m_986_io_x2 = m_294_io_cout; // @[MUL.scala 253:22]
  assign m_986_io_x3 = m_304_io_s; // @[MUL.scala 252:21]
  assign m_987_io_x1 = m_295_io_cout; // @[MUL.scala 253:22]
  assign m_987_io_x2 = m_305_io_s; // @[MUL.scala 252:21]
  assign m_987_io_x3 = m_296_io_cout; // @[MUL.scala 253:22]
  assign m_988_io_x1 = m_306_io_s; // @[MUL.scala 252:21]
  assign m_988_io_x2 = m_297_io_cout; // @[MUL.scala 253:22]
  assign m_988_io_x3 = m_307_io_s; // @[MUL.scala 252:21]
  assign m_989_io_x1 = m_298_io_cout; // @[MUL.scala 253:22]
  assign m_989_io_x2 = m_308_io_s; // @[MUL.scala 252:21]
  assign m_989_io_x3 = m_299_io_cout; // @[MUL.scala 253:22]
  assign m_990_io_x1 = m_309_io_s; // @[MUL.scala 252:21]
  assign m_990_io_x2 = m_300_io_cout; // @[MUL.scala 253:22]
  assign m_990_io_x3 = m_310_io_s; // @[MUL.scala 252:21]
  assign m_991_io_x1 = m_301_io_cout; // @[MUL.scala 253:22]
  assign m_991_io_x2 = m_311_io_s; // @[MUL.scala 252:21]
  assign m_991_io_x3 = m_302_io_cout; // @[MUL.scala 253:22]
  assign m_992_io_x1 = m_313_io_s; // @[MUL.scala 252:21]
  assign m_992_io_x2 = m_303_io_cout; // @[MUL.scala 253:22]
  assign m_992_io_x3 = m_314_io_s; // @[MUL.scala 252:21]
  assign m_993_io_x1 = m_304_io_cout; // @[MUL.scala 253:22]
  assign m_993_io_x2 = m_315_io_s; // @[MUL.scala 252:21]
  assign m_993_io_x3 = m_305_io_cout; // @[MUL.scala 253:22]
  assign m_994_io_x1 = m_316_io_s; // @[MUL.scala 252:21]
  assign m_994_io_x2 = m_306_io_cout; // @[MUL.scala 253:22]
  assign m_994_io_x3 = m_317_io_s; // @[MUL.scala 252:21]
  assign m_995_io_x1 = m_307_io_cout; // @[MUL.scala 253:22]
  assign m_995_io_x2 = m_318_io_s; // @[MUL.scala 252:21]
  assign m_995_io_x3 = m_308_io_cout; // @[MUL.scala 253:22]
  assign m_996_io_x1 = m_319_io_s; // @[MUL.scala 252:21]
  assign m_996_io_x2 = m_309_io_cout; // @[MUL.scala 253:22]
  assign m_996_io_x3 = m_320_io_s; // @[MUL.scala 252:21]
  assign m_997_io_x1 = m_310_io_cout; // @[MUL.scala 253:22]
  assign m_997_io_x2 = m_321_io_s; // @[MUL.scala 252:21]
  assign m_997_io_x3 = m_311_io_cout; // @[MUL.scala 253:22]
  assign m_998_io_in_0 = m_322_io_out_0; // @[MUL.scala 125:16]
  assign m_998_io_in_1 = m_312_io_out_1; // @[MUL.scala 126:16]
  assign m_999_io_x1 = m_323_io_s; // @[MUL.scala 252:21]
  assign m_999_io_x2 = m_313_io_cout; // @[MUL.scala 253:22]
  assign m_999_io_x3 = m_324_io_s; // @[MUL.scala 252:21]
  assign m_1000_io_x1 = m_314_io_cout; // @[MUL.scala 253:22]
  assign m_1000_io_x2 = m_325_io_s; // @[MUL.scala 252:21]
  assign m_1000_io_x3 = m_315_io_cout; // @[MUL.scala 253:22]
  assign m_1001_io_x1 = m_326_io_s; // @[MUL.scala 252:21]
  assign m_1001_io_x2 = m_316_io_cout; // @[MUL.scala 253:22]
  assign m_1001_io_x3 = m_327_io_s; // @[MUL.scala 252:21]
  assign m_1002_io_x1 = m_317_io_cout; // @[MUL.scala 253:22]
  assign m_1002_io_x2 = m_328_io_s; // @[MUL.scala 252:21]
  assign m_1002_io_x3 = m_318_io_cout; // @[MUL.scala 253:22]
  assign m_1003_io_x1 = m_329_io_s; // @[MUL.scala 252:21]
  assign m_1003_io_x2 = m_319_io_cout; // @[MUL.scala 253:22]
  assign m_1003_io_x3 = m_330_io_s; // @[MUL.scala 252:21]
  assign m_1004_io_x1 = m_320_io_cout; // @[MUL.scala 253:22]
  assign m_1004_io_x2 = m_331_io_s; // @[MUL.scala 252:21]
  assign m_1004_io_x3 = m_321_io_cout; // @[MUL.scala 253:22]
  assign m_1005_io_in_0 = m_332_io_s; // @[MUL.scala 252:21]
  assign m_1005_io_in_1 = m_322_io_out_1; // @[MUL.scala 126:16]
  assign m_1006_io_x1 = m_333_io_s; // @[MUL.scala 252:21]
  assign m_1006_io_x2 = m_323_io_cout; // @[MUL.scala 253:22]
  assign m_1006_io_x3 = m_334_io_s; // @[MUL.scala 252:21]
  assign m_1007_io_x1 = m_324_io_cout; // @[MUL.scala 253:22]
  assign m_1007_io_x2 = m_335_io_s; // @[MUL.scala 252:21]
  assign m_1007_io_x3 = m_325_io_cout; // @[MUL.scala 253:22]
  assign m_1008_io_x1 = m_336_io_s; // @[MUL.scala 252:21]
  assign m_1008_io_x2 = m_326_io_cout; // @[MUL.scala 253:22]
  assign m_1008_io_x3 = m_337_io_s; // @[MUL.scala 252:21]
  assign m_1009_io_x1 = m_327_io_cout; // @[MUL.scala 253:22]
  assign m_1009_io_x2 = m_338_io_s; // @[MUL.scala 252:21]
  assign m_1009_io_x3 = m_328_io_cout; // @[MUL.scala 253:22]
  assign m_1010_io_x1 = m_339_io_s; // @[MUL.scala 252:21]
  assign m_1010_io_x2 = m_329_io_cout; // @[MUL.scala 253:22]
  assign m_1010_io_x3 = m_340_io_s; // @[MUL.scala 252:21]
  assign m_1011_io_x1 = m_330_io_cout; // @[MUL.scala 253:22]
  assign m_1011_io_x2 = m_341_io_s; // @[MUL.scala 252:21]
  assign m_1011_io_x3 = m_331_io_cout; // @[MUL.scala 253:22]
  assign m_1012_io_in_0 = m_342_io_s; // @[MUL.scala 252:21]
  assign m_1012_io_in_1 = m_332_io_cout; // @[MUL.scala 253:22]
  assign m_1013_io_x1 = m_343_io_s; // @[MUL.scala 252:21]
  assign m_1013_io_x2 = m_333_io_cout; // @[MUL.scala 253:22]
  assign m_1013_io_x3 = m_344_io_s; // @[MUL.scala 252:21]
  assign m_1014_io_x1 = m_334_io_cout; // @[MUL.scala 253:22]
  assign m_1014_io_x2 = m_345_io_s; // @[MUL.scala 252:21]
  assign m_1014_io_x3 = m_335_io_cout; // @[MUL.scala 253:22]
  assign m_1015_io_x1 = m_346_io_s; // @[MUL.scala 252:21]
  assign m_1015_io_x2 = m_336_io_cout; // @[MUL.scala 253:22]
  assign m_1015_io_x3 = m_347_io_s; // @[MUL.scala 252:21]
  assign m_1016_io_x1 = m_337_io_cout; // @[MUL.scala 253:22]
  assign m_1016_io_x2 = m_348_io_s; // @[MUL.scala 252:21]
  assign m_1016_io_x3 = m_338_io_cout; // @[MUL.scala 253:22]
  assign m_1017_io_x1 = m_349_io_s; // @[MUL.scala 252:21]
  assign m_1017_io_x2 = m_339_io_cout; // @[MUL.scala 253:22]
  assign m_1017_io_x3 = m_350_io_s; // @[MUL.scala 252:21]
  assign m_1018_io_x1 = m_340_io_cout; // @[MUL.scala 253:22]
  assign m_1018_io_x2 = m_351_io_s; // @[MUL.scala 252:21]
  assign m_1018_io_x3 = m_341_io_cout; // @[MUL.scala 253:22]
  assign m_1019_io_x1 = m_352_io_s; // @[MUL.scala 252:21]
  assign m_1019_io_x2 = m_342_io_cout; // @[MUL.scala 253:22]
  assign m_1019_io_x3 = r_958; // @[MUL.scala 105:13]
  assign m_1020_io_x1 = m_353_io_s; // @[MUL.scala 252:21]
  assign m_1020_io_x2 = m_343_io_cout; // @[MUL.scala 253:22]
  assign m_1020_io_x3 = m_354_io_s; // @[MUL.scala 252:21]
  assign m_1021_io_x1 = m_344_io_cout; // @[MUL.scala 253:22]
  assign m_1021_io_x2 = m_355_io_s; // @[MUL.scala 252:21]
  assign m_1021_io_x3 = m_345_io_cout; // @[MUL.scala 253:22]
  assign m_1022_io_x1 = m_356_io_s; // @[MUL.scala 252:21]
  assign m_1022_io_x2 = m_346_io_cout; // @[MUL.scala 253:22]
  assign m_1022_io_x3 = m_357_io_s; // @[MUL.scala 252:21]
  assign m_1023_io_x1 = m_347_io_cout; // @[MUL.scala 253:22]
  assign m_1023_io_x2 = m_358_io_s; // @[MUL.scala 252:21]
  assign m_1023_io_x3 = m_348_io_cout; // @[MUL.scala 253:22]
  assign m_1024_io_x1 = m_359_io_s; // @[MUL.scala 252:21]
  assign m_1024_io_x2 = m_349_io_cout; // @[MUL.scala 253:22]
  assign m_1024_io_x3 = m_360_io_s; // @[MUL.scala 252:21]
  assign m_1025_io_x1 = m_350_io_cout; // @[MUL.scala 253:22]
  assign m_1025_io_x2 = m_361_io_s; // @[MUL.scala 252:21]
  assign m_1025_io_x3 = m_351_io_cout; // @[MUL.scala 253:22]
  assign m_1026_io_x1 = m_362_io_s; // @[MUL.scala 252:21]
  assign m_1026_io_x2 = m_352_io_cout; // @[MUL.scala 253:22]
  assign m_1026_io_x3 = r_989; // @[MUL.scala 105:13]
  assign m_1027_io_x1 = m_363_io_s; // @[MUL.scala 252:21]
  assign m_1027_io_x2 = m_353_io_cout; // @[MUL.scala 253:22]
  assign m_1027_io_x3 = m_364_io_s; // @[MUL.scala 252:21]
  assign m_1028_io_x1 = m_354_io_cout; // @[MUL.scala 253:22]
  assign m_1028_io_x2 = m_365_io_s; // @[MUL.scala 252:21]
  assign m_1028_io_x3 = m_355_io_cout; // @[MUL.scala 253:22]
  assign m_1029_io_x1 = m_366_io_s; // @[MUL.scala 252:21]
  assign m_1029_io_x2 = m_356_io_cout; // @[MUL.scala 253:22]
  assign m_1029_io_x3 = m_367_io_s; // @[MUL.scala 252:21]
  assign m_1030_io_x1 = m_357_io_cout; // @[MUL.scala 253:22]
  assign m_1030_io_x2 = m_368_io_s; // @[MUL.scala 252:21]
  assign m_1030_io_x3 = m_358_io_cout; // @[MUL.scala 253:22]
  assign m_1031_io_x1 = m_369_io_s; // @[MUL.scala 252:21]
  assign m_1031_io_x2 = m_359_io_cout; // @[MUL.scala 253:22]
  assign m_1031_io_x3 = m_370_io_s; // @[MUL.scala 252:21]
  assign m_1032_io_x1 = m_360_io_cout; // @[MUL.scala 253:22]
  assign m_1032_io_x2 = m_371_io_s; // @[MUL.scala 252:21]
  assign m_1032_io_x3 = m_361_io_cout; // @[MUL.scala 253:22]
  assign m_1033_io_x1 = m_372_io_s; // @[MUL.scala 252:21]
  assign m_1033_io_x2 = m_362_io_cout; // @[MUL.scala 253:22]
  assign m_1033_io_x3 = m_373_io_out_0; // @[MUL.scala 105:13]
  assign m_1034_io_x1 = m_374_io_s; // @[MUL.scala 252:21]
  assign m_1034_io_x2 = m_363_io_cout; // @[MUL.scala 253:22]
  assign m_1034_io_x3 = m_375_io_s; // @[MUL.scala 252:21]
  assign m_1035_io_x1 = m_364_io_cout; // @[MUL.scala 253:22]
  assign m_1035_io_x2 = m_376_io_s; // @[MUL.scala 252:21]
  assign m_1035_io_x3 = m_365_io_cout; // @[MUL.scala 253:22]
  assign m_1036_io_x1 = m_377_io_s; // @[MUL.scala 252:21]
  assign m_1036_io_x2 = m_366_io_cout; // @[MUL.scala 253:22]
  assign m_1036_io_x3 = m_378_io_s; // @[MUL.scala 252:21]
  assign m_1037_io_x1 = m_367_io_cout; // @[MUL.scala 253:22]
  assign m_1037_io_x2 = m_379_io_s; // @[MUL.scala 252:21]
  assign m_1037_io_x3 = m_368_io_cout; // @[MUL.scala 253:22]
  assign m_1038_io_x1 = m_380_io_s; // @[MUL.scala 252:21]
  assign m_1038_io_x2 = m_369_io_cout; // @[MUL.scala 253:22]
  assign m_1038_io_x3 = m_381_io_s; // @[MUL.scala 252:21]
  assign m_1039_io_x1 = m_370_io_cout; // @[MUL.scala 253:22]
  assign m_1039_io_x2 = m_382_io_s; // @[MUL.scala 252:21]
  assign m_1039_io_x3 = m_371_io_cout; // @[MUL.scala 253:22]
  assign m_1040_io_x1 = m_383_io_s; // @[MUL.scala 252:21]
  assign m_1040_io_x2 = m_372_io_cout; // @[MUL.scala 253:22]
  assign m_1040_io_x3 = m_384_io_out_0; // @[MUL.scala 105:13]
  assign m_1041_io_x1 = m_385_io_s; // @[MUL.scala 252:21]
  assign m_1041_io_x2 = m_374_io_cout; // @[MUL.scala 253:22]
  assign m_1041_io_x3 = m_386_io_s; // @[MUL.scala 252:21]
  assign m_1042_io_x1 = m_375_io_cout; // @[MUL.scala 253:22]
  assign m_1042_io_x2 = m_387_io_s; // @[MUL.scala 252:21]
  assign m_1042_io_x3 = m_376_io_cout; // @[MUL.scala 253:22]
  assign m_1043_io_x1 = m_388_io_s; // @[MUL.scala 252:21]
  assign m_1043_io_x2 = m_377_io_cout; // @[MUL.scala 253:22]
  assign m_1043_io_x3 = m_389_io_s; // @[MUL.scala 252:21]
  assign m_1044_io_x1 = m_378_io_cout; // @[MUL.scala 253:22]
  assign m_1044_io_x2 = m_390_io_s; // @[MUL.scala 252:21]
  assign m_1044_io_x3 = m_379_io_cout; // @[MUL.scala 253:22]
  assign m_1045_io_x1 = m_391_io_s; // @[MUL.scala 252:21]
  assign m_1045_io_x2 = m_380_io_cout; // @[MUL.scala 253:22]
  assign m_1045_io_x3 = m_392_io_s; // @[MUL.scala 252:21]
  assign m_1046_io_x1 = m_381_io_cout; // @[MUL.scala 253:22]
  assign m_1046_io_x2 = m_393_io_s; // @[MUL.scala 252:21]
  assign m_1046_io_x3 = m_382_io_cout; // @[MUL.scala 253:22]
  assign m_1047_io_x1 = m_394_io_s; // @[MUL.scala 252:21]
  assign m_1047_io_x2 = m_383_io_cout; // @[MUL.scala 253:22]
  assign m_1047_io_x3 = m_395_io_s; // @[MUL.scala 252:21]
  assign m_1048_io_x1 = m_396_io_s; // @[MUL.scala 252:21]
  assign m_1048_io_x2 = m_385_io_cout; // @[MUL.scala 253:22]
  assign m_1048_io_x3 = m_397_io_s; // @[MUL.scala 252:21]
  assign m_1049_io_x1 = m_386_io_cout; // @[MUL.scala 253:22]
  assign m_1049_io_x2 = m_398_io_s; // @[MUL.scala 252:21]
  assign m_1049_io_x3 = m_387_io_cout; // @[MUL.scala 253:22]
  assign m_1050_io_x1 = m_399_io_s; // @[MUL.scala 252:21]
  assign m_1050_io_x2 = m_388_io_cout; // @[MUL.scala 253:22]
  assign m_1050_io_x3 = m_400_io_s; // @[MUL.scala 252:21]
  assign m_1051_io_x1 = m_389_io_cout; // @[MUL.scala 253:22]
  assign m_1051_io_x2 = m_401_io_s; // @[MUL.scala 252:21]
  assign m_1051_io_x3 = m_390_io_cout; // @[MUL.scala 253:22]
  assign m_1052_io_x1 = m_402_io_s; // @[MUL.scala 252:21]
  assign m_1052_io_x2 = m_391_io_cout; // @[MUL.scala 253:22]
  assign m_1052_io_x3 = m_403_io_s; // @[MUL.scala 252:21]
  assign m_1053_io_x1 = m_392_io_cout; // @[MUL.scala 253:22]
  assign m_1053_io_x2 = m_404_io_s; // @[MUL.scala 252:21]
  assign m_1053_io_x3 = m_393_io_cout; // @[MUL.scala 253:22]
  assign m_1054_io_x1 = m_405_io_s; // @[MUL.scala 252:21]
  assign m_1054_io_x2 = m_394_io_cout; // @[MUL.scala 253:22]
  assign m_1054_io_x3 = m_406_io_s; // @[MUL.scala 252:21]
  assign m_1055_io_x1 = m_407_io_s; // @[MUL.scala 252:21]
  assign m_1055_io_x2 = m_396_io_cout; // @[MUL.scala 253:22]
  assign m_1055_io_x3 = m_408_io_s; // @[MUL.scala 252:21]
  assign m_1056_io_x1 = m_397_io_cout; // @[MUL.scala 253:22]
  assign m_1056_io_x2 = m_409_io_s; // @[MUL.scala 252:21]
  assign m_1056_io_x3 = m_398_io_cout; // @[MUL.scala 253:22]
  assign m_1057_io_x1 = m_410_io_s; // @[MUL.scala 252:21]
  assign m_1057_io_x2 = m_399_io_cout; // @[MUL.scala 253:22]
  assign m_1057_io_x3 = m_411_io_s; // @[MUL.scala 252:21]
  assign m_1058_io_x1 = m_400_io_cout; // @[MUL.scala 253:22]
  assign m_1058_io_x2 = m_412_io_s; // @[MUL.scala 252:21]
  assign m_1058_io_x3 = m_401_io_cout; // @[MUL.scala 253:22]
  assign m_1059_io_x1 = m_413_io_s; // @[MUL.scala 252:21]
  assign m_1059_io_x2 = m_402_io_cout; // @[MUL.scala 253:22]
  assign m_1059_io_x3 = m_414_io_s; // @[MUL.scala 252:21]
  assign m_1060_io_x1 = m_403_io_cout; // @[MUL.scala 253:22]
  assign m_1060_io_x2 = m_415_io_s; // @[MUL.scala 252:21]
  assign m_1060_io_x3 = m_404_io_cout; // @[MUL.scala 253:22]
  assign m_1061_io_x1 = m_416_io_s; // @[MUL.scala 252:21]
  assign m_1061_io_x2 = m_405_io_cout; // @[MUL.scala 253:22]
  assign m_1061_io_x3 = m_417_io_s; // @[MUL.scala 252:21]
  assign m_1062_io_x1 = m_418_io_s; // @[MUL.scala 252:21]
  assign m_1062_io_x2 = m_407_io_cout; // @[MUL.scala 253:22]
  assign m_1062_io_x3 = m_419_io_s; // @[MUL.scala 252:21]
  assign m_1063_io_x1 = m_408_io_cout; // @[MUL.scala 253:22]
  assign m_1063_io_x2 = m_420_io_s; // @[MUL.scala 252:21]
  assign m_1063_io_x3 = m_409_io_cout; // @[MUL.scala 253:22]
  assign m_1064_io_x1 = m_421_io_s; // @[MUL.scala 252:21]
  assign m_1064_io_x2 = m_410_io_cout; // @[MUL.scala 253:22]
  assign m_1064_io_x3 = m_422_io_s; // @[MUL.scala 252:21]
  assign m_1065_io_x1 = m_411_io_cout; // @[MUL.scala 253:22]
  assign m_1065_io_x2 = m_423_io_s; // @[MUL.scala 252:21]
  assign m_1065_io_x3 = m_412_io_cout; // @[MUL.scala 253:22]
  assign m_1066_io_x1 = m_424_io_s; // @[MUL.scala 252:21]
  assign m_1066_io_x2 = m_413_io_cout; // @[MUL.scala 253:22]
  assign m_1066_io_x3 = m_425_io_s; // @[MUL.scala 252:21]
  assign m_1067_io_x1 = m_414_io_cout; // @[MUL.scala 253:22]
  assign m_1067_io_x2 = m_426_io_s; // @[MUL.scala 252:21]
  assign m_1067_io_x3 = m_415_io_cout; // @[MUL.scala 253:22]
  assign m_1068_io_x1 = m_427_io_s; // @[MUL.scala 252:21]
  assign m_1068_io_x2 = m_416_io_cout; // @[MUL.scala 253:22]
  assign m_1068_io_x3 = m_428_io_s; // @[MUL.scala 252:21]
  assign m_1069_io_x1 = m_429_io_s; // @[MUL.scala 252:21]
  assign m_1069_io_x2 = m_418_io_cout; // @[MUL.scala 253:22]
  assign m_1069_io_x3 = m_430_io_s; // @[MUL.scala 252:21]
  assign m_1070_io_x1 = m_419_io_cout; // @[MUL.scala 253:22]
  assign m_1070_io_x2 = m_431_io_s; // @[MUL.scala 252:21]
  assign m_1070_io_x3 = m_420_io_cout; // @[MUL.scala 253:22]
  assign m_1071_io_x1 = m_432_io_s; // @[MUL.scala 252:21]
  assign m_1071_io_x2 = m_421_io_cout; // @[MUL.scala 253:22]
  assign m_1071_io_x3 = m_433_io_s; // @[MUL.scala 252:21]
  assign m_1072_io_x1 = m_422_io_cout; // @[MUL.scala 253:22]
  assign m_1072_io_x2 = m_434_io_s; // @[MUL.scala 252:21]
  assign m_1072_io_x3 = m_423_io_cout; // @[MUL.scala 253:22]
  assign m_1073_io_x1 = m_435_io_s; // @[MUL.scala 252:21]
  assign m_1073_io_x2 = m_424_io_cout; // @[MUL.scala 253:22]
  assign m_1073_io_x3 = m_436_io_s; // @[MUL.scala 252:21]
  assign m_1074_io_x1 = m_425_io_cout; // @[MUL.scala 253:22]
  assign m_1074_io_x2 = m_437_io_s; // @[MUL.scala 252:21]
  assign m_1074_io_x3 = m_426_io_cout; // @[MUL.scala 253:22]
  assign m_1075_io_x1 = m_438_io_s; // @[MUL.scala 252:21]
  assign m_1075_io_x2 = m_427_io_cout; // @[MUL.scala 253:22]
  assign m_1075_io_x3 = m_439_io_s; // @[MUL.scala 252:21]
  assign m_1076_io_x1 = m_440_io_s; // @[MUL.scala 252:21]
  assign m_1076_io_x2 = m_429_io_cout; // @[MUL.scala 253:22]
  assign m_1076_io_x3 = m_441_io_s; // @[MUL.scala 252:21]
  assign m_1077_io_x1 = m_430_io_cout; // @[MUL.scala 253:22]
  assign m_1077_io_x2 = m_442_io_s; // @[MUL.scala 252:21]
  assign m_1077_io_x3 = m_431_io_cout; // @[MUL.scala 253:22]
  assign m_1078_io_x1 = m_443_io_s; // @[MUL.scala 252:21]
  assign m_1078_io_x2 = m_432_io_cout; // @[MUL.scala 253:22]
  assign m_1078_io_x3 = m_444_io_s; // @[MUL.scala 252:21]
  assign m_1079_io_x1 = m_433_io_cout; // @[MUL.scala 253:22]
  assign m_1079_io_x2 = m_445_io_s; // @[MUL.scala 252:21]
  assign m_1079_io_x3 = m_434_io_cout; // @[MUL.scala 253:22]
  assign m_1080_io_x1 = m_446_io_s; // @[MUL.scala 252:21]
  assign m_1080_io_x2 = m_435_io_cout; // @[MUL.scala 253:22]
  assign m_1080_io_x3 = m_447_io_s; // @[MUL.scala 252:21]
  assign m_1081_io_x1 = m_436_io_cout; // @[MUL.scala 253:22]
  assign m_1081_io_x2 = m_448_io_s; // @[MUL.scala 252:21]
  assign m_1081_io_x3 = m_437_io_cout; // @[MUL.scala 253:22]
  assign m_1082_io_x1 = m_449_io_s; // @[MUL.scala 252:21]
  assign m_1082_io_x2 = m_438_io_cout; // @[MUL.scala 253:22]
  assign m_1082_io_x3 = m_450_io_s; // @[MUL.scala 252:21]
  assign m_1083_io_x1 = m_451_io_s; // @[MUL.scala 252:21]
  assign m_1083_io_x2 = m_440_io_cout; // @[MUL.scala 253:22]
  assign m_1083_io_x3 = m_452_io_s; // @[MUL.scala 252:21]
  assign m_1084_io_x1 = m_441_io_cout; // @[MUL.scala 253:22]
  assign m_1084_io_x2 = m_453_io_s; // @[MUL.scala 252:21]
  assign m_1084_io_x3 = m_442_io_cout; // @[MUL.scala 253:22]
  assign m_1085_io_x1 = m_454_io_s; // @[MUL.scala 252:21]
  assign m_1085_io_x2 = m_443_io_cout; // @[MUL.scala 253:22]
  assign m_1085_io_x3 = m_455_io_s; // @[MUL.scala 252:21]
  assign m_1086_io_x1 = m_444_io_cout; // @[MUL.scala 253:22]
  assign m_1086_io_x2 = m_456_io_s; // @[MUL.scala 252:21]
  assign m_1086_io_x3 = m_445_io_cout; // @[MUL.scala 253:22]
  assign m_1087_io_x1 = m_457_io_s; // @[MUL.scala 252:21]
  assign m_1087_io_x2 = m_446_io_cout; // @[MUL.scala 253:22]
  assign m_1087_io_x3 = m_458_io_s; // @[MUL.scala 252:21]
  assign m_1088_io_x1 = m_447_io_cout; // @[MUL.scala 253:22]
  assign m_1088_io_x2 = m_459_io_s; // @[MUL.scala 252:21]
  assign m_1088_io_x3 = m_448_io_cout; // @[MUL.scala 253:22]
  assign m_1089_io_x1 = m_460_io_s; // @[MUL.scala 252:21]
  assign m_1089_io_x2 = m_449_io_cout; // @[MUL.scala 253:22]
  assign m_1089_io_x3 = m_461_io_s; // @[MUL.scala 252:21]
  assign m_1090_io_x1 = m_462_io_s; // @[MUL.scala 252:21]
  assign m_1090_io_x2 = m_451_io_cout; // @[MUL.scala 253:22]
  assign m_1090_io_x3 = m_463_io_s; // @[MUL.scala 252:21]
  assign m_1091_io_x1 = m_452_io_cout; // @[MUL.scala 253:22]
  assign m_1091_io_x2 = m_464_io_s; // @[MUL.scala 252:21]
  assign m_1091_io_x3 = m_453_io_cout; // @[MUL.scala 253:22]
  assign m_1092_io_x1 = m_465_io_s; // @[MUL.scala 252:21]
  assign m_1092_io_x2 = m_454_io_cout; // @[MUL.scala 253:22]
  assign m_1092_io_x3 = m_466_io_s; // @[MUL.scala 252:21]
  assign m_1093_io_x1 = m_455_io_cout; // @[MUL.scala 253:22]
  assign m_1093_io_x2 = m_467_io_s; // @[MUL.scala 252:21]
  assign m_1093_io_x3 = m_456_io_cout; // @[MUL.scala 253:22]
  assign m_1094_io_x1 = m_468_io_s; // @[MUL.scala 252:21]
  assign m_1094_io_x2 = m_457_io_cout; // @[MUL.scala 253:22]
  assign m_1094_io_x3 = m_469_io_s; // @[MUL.scala 252:21]
  assign m_1095_io_x1 = m_458_io_cout; // @[MUL.scala 253:22]
  assign m_1095_io_x2 = m_470_io_s; // @[MUL.scala 252:21]
  assign m_1095_io_x3 = m_459_io_cout; // @[MUL.scala 253:22]
  assign m_1096_io_x1 = m_471_io_s; // @[MUL.scala 252:21]
  assign m_1096_io_x2 = m_460_io_cout; // @[MUL.scala 253:22]
  assign m_1096_io_x3 = m_472_io_out_0; // @[MUL.scala 105:13]
  assign m_1097_io_x1 = m_473_io_s; // @[MUL.scala 252:21]
  assign m_1097_io_x2 = m_462_io_cout; // @[MUL.scala 253:22]
  assign m_1097_io_x3 = m_474_io_s; // @[MUL.scala 252:21]
  assign m_1098_io_x1 = m_463_io_cout; // @[MUL.scala 253:22]
  assign m_1098_io_x2 = m_475_io_s; // @[MUL.scala 252:21]
  assign m_1098_io_x3 = m_464_io_cout; // @[MUL.scala 253:22]
  assign m_1099_io_x1 = m_476_io_s; // @[MUL.scala 252:21]
  assign m_1099_io_x2 = m_465_io_cout; // @[MUL.scala 253:22]
  assign m_1099_io_x3 = m_477_io_s; // @[MUL.scala 252:21]
  assign m_1100_io_x1 = m_466_io_cout; // @[MUL.scala 253:22]
  assign m_1100_io_x2 = m_478_io_s; // @[MUL.scala 252:21]
  assign m_1100_io_x3 = m_467_io_cout; // @[MUL.scala 253:22]
  assign m_1101_io_x1 = m_479_io_s; // @[MUL.scala 252:21]
  assign m_1101_io_x2 = m_468_io_cout; // @[MUL.scala 253:22]
  assign m_1101_io_x3 = m_480_io_s; // @[MUL.scala 252:21]
  assign m_1102_io_x1 = m_469_io_cout; // @[MUL.scala 253:22]
  assign m_1102_io_x2 = m_481_io_s; // @[MUL.scala 252:21]
  assign m_1102_io_x3 = m_470_io_cout; // @[MUL.scala 253:22]
  assign m_1103_io_x1 = m_482_io_s; // @[MUL.scala 252:21]
  assign m_1103_io_x2 = m_471_io_cout; // @[MUL.scala 253:22]
  assign m_1103_io_x3 = r_1347; // @[MUL.scala 105:13]
  assign m_1104_io_x1 = m_483_io_s; // @[MUL.scala 252:21]
  assign m_1104_io_x2 = m_473_io_cout; // @[MUL.scala 253:22]
  assign m_1104_io_x3 = m_484_io_s; // @[MUL.scala 252:21]
  assign m_1105_io_x1 = m_474_io_cout; // @[MUL.scala 253:22]
  assign m_1105_io_x2 = m_485_io_s; // @[MUL.scala 252:21]
  assign m_1105_io_x3 = m_475_io_cout; // @[MUL.scala 253:22]
  assign m_1106_io_x1 = m_486_io_s; // @[MUL.scala 252:21]
  assign m_1106_io_x2 = m_476_io_cout; // @[MUL.scala 253:22]
  assign m_1106_io_x3 = m_487_io_s; // @[MUL.scala 252:21]
  assign m_1107_io_x1 = m_477_io_cout; // @[MUL.scala 253:22]
  assign m_1107_io_x2 = m_488_io_s; // @[MUL.scala 252:21]
  assign m_1107_io_x3 = m_478_io_cout; // @[MUL.scala 253:22]
  assign m_1108_io_x1 = m_489_io_s; // @[MUL.scala 252:21]
  assign m_1108_io_x2 = m_479_io_cout; // @[MUL.scala 253:22]
  assign m_1108_io_x3 = m_490_io_s; // @[MUL.scala 252:21]
  assign m_1109_io_x1 = m_480_io_cout; // @[MUL.scala 253:22]
  assign m_1109_io_x2 = m_491_io_s; // @[MUL.scala 252:21]
  assign m_1109_io_x3 = m_481_io_cout; // @[MUL.scala 253:22]
  assign m_1110_io_x1 = m_492_io_s; // @[MUL.scala 252:21]
  assign m_1110_io_x2 = m_482_io_cout; // @[MUL.scala 253:22]
  assign m_1110_io_x3 = r_1378; // @[MUL.scala 105:13]
  assign m_1111_io_x1 = m_493_io_s; // @[MUL.scala 252:21]
  assign m_1111_io_x2 = m_483_io_cout; // @[MUL.scala 253:22]
  assign m_1111_io_x3 = m_494_io_s; // @[MUL.scala 252:21]
  assign m_1112_io_x1 = m_484_io_cout; // @[MUL.scala 253:22]
  assign m_1112_io_x2 = m_495_io_s; // @[MUL.scala 252:21]
  assign m_1112_io_x3 = m_485_io_cout; // @[MUL.scala 253:22]
  assign m_1113_io_x1 = m_496_io_s; // @[MUL.scala 252:21]
  assign m_1113_io_x2 = m_486_io_cout; // @[MUL.scala 253:22]
  assign m_1113_io_x3 = m_497_io_s; // @[MUL.scala 252:21]
  assign m_1114_io_x1 = m_487_io_cout; // @[MUL.scala 253:22]
  assign m_1114_io_x2 = m_498_io_s; // @[MUL.scala 252:21]
  assign m_1114_io_x3 = m_488_io_cout; // @[MUL.scala 253:22]
  assign m_1115_io_x1 = m_499_io_s; // @[MUL.scala 252:21]
  assign m_1115_io_x2 = m_489_io_cout; // @[MUL.scala 253:22]
  assign m_1115_io_x3 = m_500_io_s; // @[MUL.scala 252:21]
  assign m_1116_io_x1 = m_490_io_cout; // @[MUL.scala 253:22]
  assign m_1116_io_x2 = m_501_io_s; // @[MUL.scala 252:21]
  assign m_1116_io_x3 = m_491_io_cout; // @[MUL.scala 253:22]
  assign m_1117_io_in_0 = m_502_io_s; // @[MUL.scala 252:21]
  assign m_1117_io_in_1 = m_492_io_cout; // @[MUL.scala 253:22]
  assign m_1118_io_x1 = m_503_io_s; // @[MUL.scala 252:21]
  assign m_1118_io_x2 = m_493_io_cout; // @[MUL.scala 253:22]
  assign m_1118_io_x3 = m_504_io_s; // @[MUL.scala 252:21]
  assign m_1119_io_x1 = m_494_io_cout; // @[MUL.scala 253:22]
  assign m_1119_io_x2 = m_505_io_s; // @[MUL.scala 252:21]
  assign m_1119_io_x3 = m_495_io_cout; // @[MUL.scala 253:22]
  assign m_1120_io_x1 = m_506_io_s; // @[MUL.scala 252:21]
  assign m_1120_io_x2 = m_496_io_cout; // @[MUL.scala 253:22]
  assign m_1120_io_x3 = m_507_io_s; // @[MUL.scala 252:21]
  assign m_1121_io_x1 = m_497_io_cout; // @[MUL.scala 253:22]
  assign m_1121_io_x2 = m_508_io_s; // @[MUL.scala 252:21]
  assign m_1121_io_x3 = m_498_io_cout; // @[MUL.scala 253:22]
  assign m_1122_io_x1 = m_509_io_s; // @[MUL.scala 252:21]
  assign m_1122_io_x2 = m_499_io_cout; // @[MUL.scala 253:22]
  assign m_1122_io_x3 = m_510_io_s; // @[MUL.scala 252:21]
  assign m_1123_io_x1 = m_500_io_cout; // @[MUL.scala 253:22]
  assign m_1123_io_x2 = m_511_io_s; // @[MUL.scala 252:21]
  assign m_1123_io_x3 = m_501_io_cout; // @[MUL.scala 253:22]
  assign m_1124_io_in_0 = m_512_io_s; // @[MUL.scala 252:21]
  assign m_1124_io_in_1 = m_502_io_cout; // @[MUL.scala 253:22]
  assign m_1125_io_x1 = m_513_io_s; // @[MUL.scala 252:21]
  assign m_1125_io_x2 = m_503_io_cout; // @[MUL.scala 253:22]
  assign m_1125_io_x3 = m_514_io_s; // @[MUL.scala 252:21]
  assign m_1126_io_x1 = m_504_io_cout; // @[MUL.scala 253:22]
  assign m_1126_io_x2 = m_515_io_s; // @[MUL.scala 252:21]
  assign m_1126_io_x3 = m_505_io_cout; // @[MUL.scala 253:22]
  assign m_1127_io_x1 = m_516_io_s; // @[MUL.scala 252:21]
  assign m_1127_io_x2 = m_506_io_cout; // @[MUL.scala 253:22]
  assign m_1127_io_x3 = m_517_io_s; // @[MUL.scala 252:21]
  assign m_1128_io_x1 = m_507_io_cout; // @[MUL.scala 253:22]
  assign m_1128_io_x2 = m_518_io_s; // @[MUL.scala 252:21]
  assign m_1128_io_x3 = m_508_io_cout; // @[MUL.scala 253:22]
  assign m_1129_io_x1 = m_519_io_s; // @[MUL.scala 252:21]
  assign m_1129_io_x2 = m_509_io_cout; // @[MUL.scala 253:22]
  assign m_1129_io_x3 = m_520_io_s; // @[MUL.scala 252:21]
  assign m_1130_io_x1 = m_510_io_cout; // @[MUL.scala 253:22]
  assign m_1130_io_x2 = m_521_io_s; // @[MUL.scala 252:21]
  assign m_1130_io_x3 = m_511_io_cout; // @[MUL.scala 253:22]
  assign m_1131_io_in_0 = m_522_io_out_0; // @[MUL.scala 125:16]
  assign m_1131_io_in_1 = m_512_io_cout; // @[MUL.scala 253:22]
  assign m_1132_io_x1 = m_523_io_s; // @[MUL.scala 252:21]
  assign m_1132_io_x2 = m_513_io_cout; // @[MUL.scala 253:22]
  assign m_1132_io_x3 = m_524_io_s; // @[MUL.scala 252:21]
  assign m_1133_io_x1 = m_514_io_cout; // @[MUL.scala 253:22]
  assign m_1133_io_x2 = m_525_io_s; // @[MUL.scala 252:21]
  assign m_1133_io_x3 = m_515_io_cout; // @[MUL.scala 253:22]
  assign m_1134_io_x1 = m_526_io_s; // @[MUL.scala 252:21]
  assign m_1134_io_x2 = m_516_io_cout; // @[MUL.scala 253:22]
  assign m_1134_io_x3 = m_527_io_s; // @[MUL.scala 252:21]
  assign m_1135_io_x1 = m_517_io_cout; // @[MUL.scala 253:22]
  assign m_1135_io_x2 = m_528_io_s; // @[MUL.scala 252:21]
  assign m_1135_io_x3 = m_518_io_cout; // @[MUL.scala 253:22]
  assign m_1136_io_x1 = m_529_io_s; // @[MUL.scala 252:21]
  assign m_1136_io_x2 = m_519_io_cout; // @[MUL.scala 253:22]
  assign m_1136_io_x3 = m_530_io_s; // @[MUL.scala 252:21]
  assign m_1137_io_x1 = m_520_io_cout; // @[MUL.scala 253:22]
  assign m_1137_io_x2 = m_531_io_s; // @[MUL.scala 252:21]
  assign m_1137_io_x3 = m_521_io_cout; // @[MUL.scala 253:22]
  assign m_1138_io_in_0 = m_532_io_out_0; // @[MUL.scala 125:16]
  assign m_1138_io_in_1 = m_522_io_out_1; // @[MUL.scala 126:16]
  assign m_1139_io_x1 = m_533_io_s; // @[MUL.scala 252:21]
  assign m_1139_io_x2 = m_523_io_cout; // @[MUL.scala 253:22]
  assign m_1139_io_x3 = m_534_io_s; // @[MUL.scala 252:21]
  assign m_1140_io_x1 = m_524_io_cout; // @[MUL.scala 253:22]
  assign m_1140_io_x2 = m_535_io_s; // @[MUL.scala 252:21]
  assign m_1140_io_x3 = m_525_io_cout; // @[MUL.scala 253:22]
  assign m_1141_io_x1 = m_536_io_s; // @[MUL.scala 252:21]
  assign m_1141_io_x2 = m_526_io_cout; // @[MUL.scala 253:22]
  assign m_1141_io_x3 = m_537_io_s; // @[MUL.scala 252:21]
  assign m_1142_io_x1 = m_527_io_cout; // @[MUL.scala 253:22]
  assign m_1142_io_x2 = m_538_io_s; // @[MUL.scala 252:21]
  assign m_1142_io_x3 = m_528_io_cout; // @[MUL.scala 253:22]
  assign m_1143_io_x1 = m_539_io_s; // @[MUL.scala 252:21]
  assign m_1143_io_x2 = m_529_io_cout; // @[MUL.scala 253:22]
  assign m_1143_io_x3 = m_540_io_s; // @[MUL.scala 252:21]
  assign m_1144_io_x1 = m_530_io_cout; // @[MUL.scala 253:22]
  assign m_1144_io_x2 = m_541_io_s; // @[MUL.scala 252:21]
  assign m_1144_io_x3 = m_531_io_cout; // @[MUL.scala 253:22]
  assign m_1145_io_in_0 = r_1524; // @[MUL.scala 125:16]
  assign m_1145_io_in_1 = m_532_io_out_1; // @[MUL.scala 126:16]
  assign m_1146_io_x1 = m_542_io_s; // @[MUL.scala 252:21]
  assign m_1146_io_x2 = m_533_io_cout; // @[MUL.scala 253:22]
  assign m_1146_io_x3 = m_543_io_s; // @[MUL.scala 252:21]
  assign m_1147_io_x1 = m_534_io_cout; // @[MUL.scala 253:22]
  assign m_1147_io_x2 = m_544_io_s; // @[MUL.scala 252:21]
  assign m_1147_io_x3 = m_535_io_cout; // @[MUL.scala 253:22]
  assign m_1148_io_x1 = m_545_io_s; // @[MUL.scala 252:21]
  assign m_1148_io_x2 = m_536_io_cout; // @[MUL.scala 253:22]
  assign m_1148_io_x3 = m_546_io_s; // @[MUL.scala 252:21]
  assign m_1149_io_x1 = m_537_io_cout; // @[MUL.scala 253:22]
  assign m_1149_io_x2 = m_547_io_s; // @[MUL.scala 252:21]
  assign m_1149_io_x3 = m_538_io_cout; // @[MUL.scala 253:22]
  assign m_1150_io_x1 = m_548_io_s; // @[MUL.scala 252:21]
  assign m_1150_io_x2 = m_539_io_cout; // @[MUL.scala 253:22]
  assign m_1150_io_x3 = m_549_io_s; // @[MUL.scala 252:21]
  assign m_1151_io_x1 = m_540_io_cout; // @[MUL.scala 253:22]
  assign m_1151_io_x2 = m_550_io_s; // @[MUL.scala 252:21]
  assign m_1151_io_x3 = m_541_io_cout; // @[MUL.scala 253:22]
  assign m_1152_io_x1 = m_551_io_s; // @[MUL.scala 252:21]
  assign m_1152_io_x2 = m_542_io_cout; // @[MUL.scala 253:22]
  assign m_1152_io_x3 = m_552_io_s; // @[MUL.scala 252:21]
  assign m_1153_io_x1 = m_543_io_cout; // @[MUL.scala 253:22]
  assign m_1153_io_x2 = m_553_io_s; // @[MUL.scala 252:21]
  assign m_1153_io_x3 = m_544_io_cout; // @[MUL.scala 253:22]
  assign m_1154_io_x1 = m_554_io_s; // @[MUL.scala 252:21]
  assign m_1154_io_x2 = m_545_io_cout; // @[MUL.scala 253:22]
  assign m_1154_io_x3 = m_555_io_s; // @[MUL.scala 252:21]
  assign m_1155_io_x1 = m_546_io_cout; // @[MUL.scala 253:22]
  assign m_1155_io_x2 = m_556_io_s; // @[MUL.scala 252:21]
  assign m_1155_io_x3 = m_547_io_cout; // @[MUL.scala 253:22]
  assign m_1156_io_x1 = m_557_io_s; // @[MUL.scala 252:21]
  assign m_1156_io_x2 = m_548_io_cout; // @[MUL.scala 253:22]
  assign m_1156_io_x3 = m_558_io_s; // @[MUL.scala 252:21]
  assign m_1157_io_x1 = m_549_io_cout; // @[MUL.scala 253:22]
  assign m_1157_io_x2 = m_559_io_s; // @[MUL.scala 252:21]
  assign m_1157_io_x3 = m_550_io_cout; // @[MUL.scala 253:22]
  assign m_1158_io_x1 = m_560_io_s; // @[MUL.scala 252:21]
  assign m_1158_io_x2 = m_551_io_cout; // @[MUL.scala 253:22]
  assign m_1158_io_x3 = m_561_io_s; // @[MUL.scala 252:21]
  assign m_1159_io_x1 = m_552_io_cout; // @[MUL.scala 253:22]
  assign m_1159_io_x2 = m_562_io_s; // @[MUL.scala 252:21]
  assign m_1159_io_x3 = m_553_io_cout; // @[MUL.scala 253:22]
  assign m_1160_io_x1 = m_563_io_s; // @[MUL.scala 252:21]
  assign m_1160_io_x2 = m_554_io_cout; // @[MUL.scala 253:22]
  assign m_1160_io_x3 = m_564_io_s; // @[MUL.scala 252:21]
  assign m_1161_io_x1 = m_555_io_cout; // @[MUL.scala 253:22]
  assign m_1161_io_x2 = m_565_io_s; // @[MUL.scala 252:21]
  assign m_1161_io_x3 = m_556_io_cout; // @[MUL.scala 253:22]
  assign m_1162_io_x1 = m_566_io_s; // @[MUL.scala 252:21]
  assign m_1162_io_x2 = m_557_io_cout; // @[MUL.scala 253:22]
  assign m_1162_io_x3 = m_567_io_s; // @[MUL.scala 252:21]
  assign m_1163_io_x1 = m_558_io_cout; // @[MUL.scala 253:22]
  assign m_1163_io_x2 = m_568_io_s; // @[MUL.scala 252:21]
  assign m_1163_io_x3 = m_559_io_cout; // @[MUL.scala 253:22]
  assign m_1164_io_x1 = m_569_io_s; // @[MUL.scala 252:21]
  assign m_1164_io_x2 = m_560_io_cout; // @[MUL.scala 253:22]
  assign m_1164_io_x3 = m_570_io_s; // @[MUL.scala 252:21]
  assign m_1165_io_x1 = m_561_io_cout; // @[MUL.scala 253:22]
  assign m_1165_io_x2 = m_571_io_s; // @[MUL.scala 252:21]
  assign m_1165_io_x3 = m_562_io_cout; // @[MUL.scala 253:22]
  assign m_1166_io_x1 = m_572_io_s; // @[MUL.scala 252:21]
  assign m_1166_io_x2 = m_563_io_cout; // @[MUL.scala 253:22]
  assign m_1166_io_x3 = m_573_io_s; // @[MUL.scala 252:21]
  assign m_1167_io_x1 = m_564_io_cout; // @[MUL.scala 253:22]
  assign m_1167_io_x2 = m_574_io_s; // @[MUL.scala 252:21]
  assign m_1167_io_x3 = m_565_io_cout; // @[MUL.scala 253:22]
  assign m_1168_io_x1 = m_575_io_s; // @[MUL.scala 252:21]
  assign m_1168_io_x2 = m_566_io_cout; // @[MUL.scala 253:22]
  assign m_1168_io_x3 = m_576_io_s; // @[MUL.scala 252:21]
  assign m_1169_io_x1 = m_567_io_cout; // @[MUL.scala 253:22]
  assign m_1169_io_x2 = m_577_io_out_0; // @[MUL.scala 104:13]
  assign m_1169_io_x3 = m_568_io_cout; // @[MUL.scala 253:22]
  assign m_1170_io_x1 = m_578_io_s; // @[MUL.scala 252:21]
  assign m_1170_io_x2 = m_569_io_cout; // @[MUL.scala 253:22]
  assign m_1170_io_x3 = m_579_io_s; // @[MUL.scala 252:21]
  assign m_1171_io_x1 = m_570_io_cout; // @[MUL.scala 253:22]
  assign m_1171_io_x2 = m_580_io_s; // @[MUL.scala 252:21]
  assign m_1171_io_x3 = m_571_io_cout; // @[MUL.scala 253:22]
  assign m_1172_io_x1 = m_581_io_s; // @[MUL.scala 252:21]
  assign m_1172_io_x2 = m_572_io_cout; // @[MUL.scala 253:22]
  assign m_1172_io_x3 = m_582_io_s; // @[MUL.scala 252:21]
  assign m_1173_io_x1 = m_573_io_cout; // @[MUL.scala 253:22]
  assign m_1173_io_x2 = m_583_io_s; // @[MUL.scala 252:21]
  assign m_1173_io_x3 = m_574_io_cout; // @[MUL.scala 253:22]
  assign m_1174_io_x1 = m_584_io_s; // @[MUL.scala 252:21]
  assign m_1174_io_x2 = m_575_io_cout; // @[MUL.scala 253:22]
  assign m_1174_io_x3 = m_585_io_s; // @[MUL.scala 252:21]
  assign m_1175_io_x1 = m_576_io_cout; // @[MUL.scala 253:22]
  assign m_1175_io_x2 = m_586_io_out_0; // @[MUL.scala 104:13]
  assign m_1175_io_x3 = m_577_io_out_1; // @[MUL.scala 105:13]
  assign m_1176_io_x1 = m_587_io_s; // @[MUL.scala 252:21]
  assign m_1176_io_x2 = m_578_io_cout; // @[MUL.scala 253:22]
  assign m_1176_io_x3 = m_588_io_s; // @[MUL.scala 252:21]
  assign m_1177_io_x1 = m_579_io_cout; // @[MUL.scala 253:22]
  assign m_1177_io_x2 = m_589_io_s; // @[MUL.scala 252:21]
  assign m_1177_io_x3 = m_580_io_cout; // @[MUL.scala 253:22]
  assign m_1178_io_x1 = m_590_io_s; // @[MUL.scala 252:21]
  assign m_1178_io_x2 = m_581_io_cout; // @[MUL.scala 253:22]
  assign m_1178_io_x3 = m_591_io_s; // @[MUL.scala 252:21]
  assign m_1179_io_x1 = m_582_io_cout; // @[MUL.scala 253:22]
  assign m_1179_io_x2 = m_592_io_s; // @[MUL.scala 252:21]
  assign m_1179_io_x3 = m_583_io_cout; // @[MUL.scala 253:22]
  assign m_1180_io_x1 = m_593_io_s; // @[MUL.scala 252:21]
  assign m_1180_io_x2 = m_584_io_cout; // @[MUL.scala 253:22]
  assign m_1180_io_x3 = m_594_io_s; // @[MUL.scala 252:21]
  assign m_1181_io_x1 = m_585_io_cout; // @[MUL.scala 253:22]
  assign m_1181_io_x2 = r_1683; // @[MUL.scala 104:13]
  assign m_1181_io_x3 = m_586_io_out_1; // @[MUL.scala 105:13]
  assign m_1182_io_x1 = m_595_io_s; // @[MUL.scala 252:21]
  assign m_1182_io_x2 = m_587_io_cout; // @[MUL.scala 253:22]
  assign m_1182_io_x3 = m_596_io_s; // @[MUL.scala 252:21]
  assign m_1183_io_x1 = m_588_io_cout; // @[MUL.scala 253:22]
  assign m_1183_io_x2 = m_597_io_s; // @[MUL.scala 252:21]
  assign m_1183_io_x3 = m_589_io_cout; // @[MUL.scala 253:22]
  assign m_1184_io_x1 = m_598_io_s; // @[MUL.scala 252:21]
  assign m_1184_io_x2 = m_590_io_cout; // @[MUL.scala 253:22]
  assign m_1184_io_x3 = m_599_io_s; // @[MUL.scala 252:21]
  assign m_1185_io_x1 = m_591_io_cout; // @[MUL.scala 253:22]
  assign m_1185_io_x2 = m_600_io_s; // @[MUL.scala 252:21]
  assign m_1185_io_x3 = m_592_io_cout; // @[MUL.scala 253:22]
  assign m_1186_io_x1 = m_601_io_s; // @[MUL.scala 252:21]
  assign m_1186_io_x2 = m_593_io_cout; // @[MUL.scala 253:22]
  assign m_1186_io_x3 = m_602_io_s; // @[MUL.scala 252:21]
  assign m_1187_io_in_0 = m_594_io_cout; // @[MUL.scala 253:22]
  assign m_1187_io_in_1 = r_1708; // @[MUL.scala 126:16]
  assign m_1188_io_x1 = m_603_io_s; // @[MUL.scala 252:21]
  assign m_1188_io_x2 = m_595_io_cout; // @[MUL.scala 253:22]
  assign m_1188_io_x3 = m_604_io_s; // @[MUL.scala 252:21]
  assign m_1189_io_x1 = m_596_io_cout; // @[MUL.scala 253:22]
  assign m_1189_io_x2 = m_605_io_s; // @[MUL.scala 252:21]
  assign m_1189_io_x3 = m_597_io_cout; // @[MUL.scala 253:22]
  assign m_1190_io_x1 = m_606_io_s; // @[MUL.scala 252:21]
  assign m_1190_io_x2 = m_598_io_cout; // @[MUL.scala 253:22]
  assign m_1190_io_x3 = m_607_io_s; // @[MUL.scala 252:21]
  assign m_1191_io_x1 = m_599_io_cout; // @[MUL.scala 253:22]
  assign m_1191_io_x2 = m_608_io_s; // @[MUL.scala 252:21]
  assign m_1191_io_x3 = m_600_io_cout; // @[MUL.scala 253:22]
  assign m_1192_io_x1 = m_609_io_s; // @[MUL.scala 252:21]
  assign m_1192_io_x2 = m_601_io_cout; // @[MUL.scala 253:22]
  assign m_1192_io_x3 = m_610_io_s; // @[MUL.scala 252:21]
  assign m_1193_io_x1 = m_611_io_s; // @[MUL.scala 252:21]
  assign m_1193_io_x2 = m_603_io_cout; // @[MUL.scala 253:22]
  assign m_1193_io_x3 = m_612_io_s; // @[MUL.scala 252:21]
  assign m_1194_io_x1 = m_604_io_cout; // @[MUL.scala 253:22]
  assign m_1194_io_x2 = m_613_io_s; // @[MUL.scala 252:21]
  assign m_1194_io_x3 = m_605_io_cout; // @[MUL.scala 253:22]
  assign m_1195_io_x1 = m_614_io_s; // @[MUL.scala 252:21]
  assign m_1195_io_x2 = m_606_io_cout; // @[MUL.scala 253:22]
  assign m_1195_io_x3 = m_615_io_s; // @[MUL.scala 252:21]
  assign m_1196_io_x1 = m_607_io_cout; // @[MUL.scala 253:22]
  assign m_1196_io_x2 = m_616_io_s; // @[MUL.scala 252:21]
  assign m_1196_io_x3 = m_608_io_cout; // @[MUL.scala 253:22]
  assign m_1197_io_x1 = m_617_io_s; // @[MUL.scala 252:21]
  assign m_1197_io_x2 = m_609_io_cout; // @[MUL.scala 253:22]
  assign m_1197_io_x3 = m_618_io_s; // @[MUL.scala 252:21]
  assign m_1198_io_x1 = m_619_io_s; // @[MUL.scala 252:21]
  assign m_1198_io_x2 = m_611_io_cout; // @[MUL.scala 253:22]
  assign m_1198_io_x3 = m_620_io_s; // @[MUL.scala 252:21]
  assign m_1199_io_x1 = m_612_io_cout; // @[MUL.scala 253:22]
  assign m_1199_io_x2 = m_621_io_s; // @[MUL.scala 252:21]
  assign m_1199_io_x3 = m_613_io_cout; // @[MUL.scala 253:22]
  assign m_1200_io_x1 = m_622_io_s; // @[MUL.scala 252:21]
  assign m_1200_io_x2 = m_614_io_cout; // @[MUL.scala 253:22]
  assign m_1200_io_x3 = m_623_io_s; // @[MUL.scala 252:21]
  assign m_1201_io_x1 = m_615_io_cout; // @[MUL.scala 253:22]
  assign m_1201_io_x2 = m_624_io_s; // @[MUL.scala 252:21]
  assign m_1201_io_x3 = m_616_io_cout; // @[MUL.scala 253:22]
  assign m_1202_io_x1 = m_625_io_s; // @[MUL.scala 252:21]
  assign m_1202_io_x2 = m_617_io_cout; // @[MUL.scala 253:22]
  assign m_1202_io_x3 = m_626_io_out_0; // @[MUL.scala 105:13]
  assign m_1203_io_x1 = m_627_io_s; // @[MUL.scala 252:21]
  assign m_1203_io_x2 = m_619_io_cout; // @[MUL.scala 253:22]
  assign m_1203_io_x3 = m_628_io_s; // @[MUL.scala 252:21]
  assign m_1204_io_x1 = m_620_io_cout; // @[MUL.scala 253:22]
  assign m_1204_io_x2 = m_629_io_s; // @[MUL.scala 252:21]
  assign m_1204_io_x3 = m_621_io_cout; // @[MUL.scala 253:22]
  assign m_1205_io_x1 = m_630_io_s; // @[MUL.scala 252:21]
  assign m_1205_io_x2 = m_622_io_cout; // @[MUL.scala 253:22]
  assign m_1205_io_x3 = m_631_io_s; // @[MUL.scala 252:21]
  assign m_1206_io_x1 = m_623_io_cout; // @[MUL.scala 253:22]
  assign m_1206_io_x2 = m_632_io_s; // @[MUL.scala 252:21]
  assign m_1206_io_x3 = m_624_io_cout; // @[MUL.scala 253:22]
  assign m_1207_io_x1 = m_633_io_s; // @[MUL.scala 252:21]
  assign m_1207_io_x2 = m_625_io_cout; // @[MUL.scala 253:22]
  assign m_1207_io_x3 = m_634_io_out_0; // @[MUL.scala 105:13]
  assign m_1208_io_x1 = m_635_io_s; // @[MUL.scala 252:21]
  assign m_1208_io_x2 = m_627_io_cout; // @[MUL.scala 253:22]
  assign m_1208_io_x3 = m_636_io_s; // @[MUL.scala 252:21]
  assign m_1209_io_x1 = m_628_io_cout; // @[MUL.scala 253:22]
  assign m_1209_io_x2 = m_637_io_s; // @[MUL.scala 252:21]
  assign m_1209_io_x3 = m_629_io_cout; // @[MUL.scala 253:22]
  assign m_1210_io_x1 = m_638_io_s; // @[MUL.scala 252:21]
  assign m_1210_io_x2 = m_630_io_cout; // @[MUL.scala 253:22]
  assign m_1210_io_x3 = m_639_io_s; // @[MUL.scala 252:21]
  assign m_1211_io_x1 = m_631_io_cout; // @[MUL.scala 253:22]
  assign m_1211_io_x2 = m_640_io_s; // @[MUL.scala 252:21]
  assign m_1211_io_x3 = m_632_io_cout; // @[MUL.scala 253:22]
  assign m_1212_io_x1 = m_641_io_s; // @[MUL.scala 252:21]
  assign m_1212_io_x2 = m_633_io_cout; // @[MUL.scala 253:22]
  assign m_1212_io_x3 = r_1824; // @[MUL.scala 105:13]
  assign m_1213_io_x1 = m_642_io_s; // @[MUL.scala 252:21]
  assign m_1213_io_x2 = m_635_io_cout; // @[MUL.scala 253:22]
  assign m_1213_io_x3 = m_643_io_s; // @[MUL.scala 252:21]
  assign m_1214_io_x1 = m_636_io_cout; // @[MUL.scala 253:22]
  assign m_1214_io_x2 = m_644_io_s; // @[MUL.scala 252:21]
  assign m_1214_io_x3 = m_637_io_cout; // @[MUL.scala 253:22]
  assign m_1215_io_x1 = m_645_io_s; // @[MUL.scala 252:21]
  assign m_1215_io_x2 = m_638_io_cout; // @[MUL.scala 253:22]
  assign m_1215_io_x3 = m_646_io_s; // @[MUL.scala 252:21]
  assign m_1216_io_x1 = m_639_io_cout; // @[MUL.scala 253:22]
  assign m_1216_io_x2 = m_647_io_s; // @[MUL.scala 252:21]
  assign m_1216_io_x3 = m_640_io_cout; // @[MUL.scala 253:22]
  assign m_1217_io_x1 = m_648_io_s; // @[MUL.scala 252:21]
  assign m_1217_io_x2 = m_641_io_cout; // @[MUL.scala 253:22]
  assign m_1217_io_x3 = r_1846; // @[MUL.scala 105:13]
  assign m_1218_io_x1 = m_649_io_s; // @[MUL.scala 252:21]
  assign m_1218_io_x2 = m_642_io_cout; // @[MUL.scala 253:22]
  assign m_1218_io_x3 = m_650_io_s; // @[MUL.scala 252:21]
  assign m_1219_io_x1 = m_643_io_cout; // @[MUL.scala 253:22]
  assign m_1219_io_x2 = m_651_io_s; // @[MUL.scala 252:21]
  assign m_1219_io_x3 = m_644_io_cout; // @[MUL.scala 253:22]
  assign m_1220_io_x1 = m_652_io_s; // @[MUL.scala 252:21]
  assign m_1220_io_x2 = m_645_io_cout; // @[MUL.scala 253:22]
  assign m_1220_io_x3 = m_653_io_s; // @[MUL.scala 252:21]
  assign m_1221_io_x1 = m_646_io_cout; // @[MUL.scala 253:22]
  assign m_1221_io_x2 = m_654_io_s; // @[MUL.scala 252:21]
  assign m_1221_io_x3 = m_647_io_cout; // @[MUL.scala 253:22]
  assign m_1222_io_in_0 = m_655_io_s; // @[MUL.scala 252:21]
  assign m_1222_io_in_1 = m_648_io_cout; // @[MUL.scala 253:22]
  assign m_1223_io_x1 = m_656_io_s; // @[MUL.scala 252:21]
  assign m_1223_io_x2 = m_649_io_cout; // @[MUL.scala 253:22]
  assign m_1223_io_x3 = m_657_io_s; // @[MUL.scala 252:21]
  assign m_1224_io_x1 = m_650_io_cout; // @[MUL.scala 253:22]
  assign m_1224_io_x2 = m_658_io_s; // @[MUL.scala 252:21]
  assign m_1224_io_x3 = m_651_io_cout; // @[MUL.scala 253:22]
  assign m_1225_io_x1 = m_659_io_s; // @[MUL.scala 252:21]
  assign m_1225_io_x2 = m_652_io_cout; // @[MUL.scala 253:22]
  assign m_1225_io_x3 = m_660_io_s; // @[MUL.scala 252:21]
  assign m_1226_io_x1 = m_653_io_cout; // @[MUL.scala 253:22]
  assign m_1226_io_x2 = m_661_io_s; // @[MUL.scala 252:21]
  assign m_1226_io_x3 = m_654_io_cout; // @[MUL.scala 253:22]
  assign m_1227_io_in_0 = m_662_io_s; // @[MUL.scala 252:21]
  assign m_1227_io_in_1 = m_655_io_cout; // @[MUL.scala 253:22]
  assign m_1228_io_x1 = m_663_io_s; // @[MUL.scala 252:21]
  assign m_1228_io_x2 = m_656_io_cout; // @[MUL.scala 253:22]
  assign m_1228_io_x3 = m_664_io_s; // @[MUL.scala 252:21]
  assign m_1229_io_x1 = m_657_io_cout; // @[MUL.scala 253:22]
  assign m_1229_io_x2 = m_665_io_s; // @[MUL.scala 252:21]
  assign m_1229_io_x3 = m_658_io_cout; // @[MUL.scala 253:22]
  assign m_1230_io_x1 = m_666_io_s; // @[MUL.scala 252:21]
  assign m_1230_io_x2 = m_659_io_cout; // @[MUL.scala 253:22]
  assign m_1230_io_x3 = m_667_io_s; // @[MUL.scala 252:21]
  assign m_1231_io_x1 = m_660_io_cout; // @[MUL.scala 253:22]
  assign m_1231_io_x2 = m_668_io_s; // @[MUL.scala 252:21]
  assign m_1231_io_x3 = m_661_io_cout; // @[MUL.scala 253:22]
  assign m_1232_io_in_0 = m_669_io_out_0; // @[MUL.scala 125:16]
  assign m_1232_io_in_1 = m_662_io_cout; // @[MUL.scala 253:22]
  assign m_1233_io_x1 = m_670_io_s; // @[MUL.scala 252:21]
  assign m_1233_io_x2 = m_663_io_cout; // @[MUL.scala 253:22]
  assign m_1233_io_x3 = m_671_io_s; // @[MUL.scala 252:21]
  assign m_1234_io_x1 = m_664_io_cout; // @[MUL.scala 253:22]
  assign m_1234_io_x2 = m_672_io_s; // @[MUL.scala 252:21]
  assign m_1234_io_x3 = m_665_io_cout; // @[MUL.scala 253:22]
  assign m_1235_io_x1 = m_673_io_s; // @[MUL.scala 252:21]
  assign m_1235_io_x2 = m_666_io_cout; // @[MUL.scala 253:22]
  assign m_1235_io_x3 = m_674_io_s; // @[MUL.scala 252:21]
  assign m_1236_io_x1 = m_667_io_cout; // @[MUL.scala 253:22]
  assign m_1236_io_x2 = m_675_io_s; // @[MUL.scala 252:21]
  assign m_1236_io_x3 = m_668_io_cout; // @[MUL.scala 253:22]
  assign m_1237_io_in_0 = m_676_io_out_0; // @[MUL.scala 125:16]
  assign m_1237_io_in_1 = m_669_io_out_1; // @[MUL.scala 126:16]
  assign m_1238_io_x1 = m_677_io_s; // @[MUL.scala 252:21]
  assign m_1238_io_x2 = m_670_io_cout; // @[MUL.scala 253:22]
  assign m_1238_io_x3 = m_678_io_s; // @[MUL.scala 252:21]
  assign m_1239_io_x1 = m_671_io_cout; // @[MUL.scala 253:22]
  assign m_1239_io_x2 = m_679_io_s; // @[MUL.scala 252:21]
  assign m_1239_io_x3 = m_672_io_cout; // @[MUL.scala 253:22]
  assign m_1240_io_x1 = m_680_io_s; // @[MUL.scala 252:21]
  assign m_1240_io_x2 = m_673_io_cout; // @[MUL.scala 253:22]
  assign m_1240_io_x3 = m_681_io_s; // @[MUL.scala 252:21]
  assign m_1241_io_x1 = m_674_io_cout; // @[MUL.scala 253:22]
  assign m_1241_io_x2 = m_682_io_s; // @[MUL.scala 252:21]
  assign m_1241_io_x3 = m_675_io_cout; // @[MUL.scala 253:22]
  assign m_1242_io_in_0 = r_1947; // @[MUL.scala 125:16]
  assign m_1242_io_in_1 = m_676_io_out_1; // @[MUL.scala 126:16]
  assign m_1243_io_x1 = m_683_io_s; // @[MUL.scala 252:21]
  assign m_1243_io_x2 = m_677_io_cout; // @[MUL.scala 253:22]
  assign m_1243_io_x3 = m_684_io_s; // @[MUL.scala 252:21]
  assign m_1244_io_x1 = m_678_io_cout; // @[MUL.scala 253:22]
  assign m_1244_io_x2 = m_685_io_s; // @[MUL.scala 252:21]
  assign m_1244_io_x3 = m_679_io_cout; // @[MUL.scala 253:22]
  assign m_1245_io_x1 = m_686_io_s; // @[MUL.scala 252:21]
  assign m_1245_io_x2 = m_680_io_cout; // @[MUL.scala 253:22]
  assign m_1245_io_x3 = m_687_io_s; // @[MUL.scala 252:21]
  assign m_1246_io_x1 = m_681_io_cout; // @[MUL.scala 253:22]
  assign m_1246_io_x2 = m_688_io_s; // @[MUL.scala 252:21]
  assign m_1246_io_x3 = m_682_io_cout; // @[MUL.scala 253:22]
  assign m_1247_io_x1 = m_689_io_s; // @[MUL.scala 252:21]
  assign m_1247_io_x2 = m_683_io_cout; // @[MUL.scala 253:22]
  assign m_1247_io_x3 = m_690_io_s; // @[MUL.scala 252:21]
  assign m_1248_io_x1 = m_684_io_cout; // @[MUL.scala 253:22]
  assign m_1248_io_x2 = m_691_io_s; // @[MUL.scala 252:21]
  assign m_1248_io_x3 = m_685_io_cout; // @[MUL.scala 253:22]
  assign m_1249_io_x1 = m_692_io_s; // @[MUL.scala 252:21]
  assign m_1249_io_x2 = m_686_io_cout; // @[MUL.scala 253:22]
  assign m_1249_io_x3 = m_693_io_s; // @[MUL.scala 252:21]
  assign m_1250_io_x1 = m_687_io_cout; // @[MUL.scala 253:22]
  assign m_1250_io_x2 = m_694_io_s; // @[MUL.scala 252:21]
  assign m_1250_io_x3 = m_688_io_cout; // @[MUL.scala 253:22]
  assign m_1251_io_x1 = m_695_io_s; // @[MUL.scala 252:21]
  assign m_1251_io_x2 = m_689_io_cout; // @[MUL.scala 253:22]
  assign m_1251_io_x3 = m_696_io_s; // @[MUL.scala 252:21]
  assign m_1252_io_x1 = m_690_io_cout; // @[MUL.scala 253:22]
  assign m_1252_io_x2 = m_697_io_s; // @[MUL.scala 252:21]
  assign m_1252_io_x3 = m_691_io_cout; // @[MUL.scala 253:22]
  assign m_1253_io_x1 = m_698_io_s; // @[MUL.scala 252:21]
  assign m_1253_io_x2 = m_692_io_cout; // @[MUL.scala 253:22]
  assign m_1253_io_x3 = m_699_io_s; // @[MUL.scala 252:21]
  assign m_1254_io_x1 = m_693_io_cout; // @[MUL.scala 253:22]
  assign m_1254_io_x2 = m_700_io_s; // @[MUL.scala 252:21]
  assign m_1254_io_x3 = m_694_io_cout; // @[MUL.scala 253:22]
  assign m_1255_io_x1 = m_701_io_s; // @[MUL.scala 252:21]
  assign m_1255_io_x2 = m_695_io_cout; // @[MUL.scala 253:22]
  assign m_1255_io_x3 = m_702_io_s; // @[MUL.scala 252:21]
  assign m_1256_io_x1 = m_696_io_cout; // @[MUL.scala 253:22]
  assign m_1256_io_x2 = m_703_io_s; // @[MUL.scala 252:21]
  assign m_1256_io_x3 = m_697_io_cout; // @[MUL.scala 253:22]
  assign m_1257_io_x1 = m_704_io_s; // @[MUL.scala 252:21]
  assign m_1257_io_x2 = m_698_io_cout; // @[MUL.scala 253:22]
  assign m_1257_io_x3 = m_705_io_s; // @[MUL.scala 252:21]
  assign m_1258_io_x1 = m_699_io_cout; // @[MUL.scala 253:22]
  assign m_1258_io_x2 = m_706_io_out_0; // @[MUL.scala 104:13]
  assign m_1258_io_x3 = m_700_io_cout; // @[MUL.scala 253:22]
  assign m_1259_io_x1 = m_707_io_s; // @[MUL.scala 252:21]
  assign m_1259_io_x2 = m_701_io_cout; // @[MUL.scala 253:22]
  assign m_1259_io_x3 = m_708_io_s; // @[MUL.scala 252:21]
  assign m_1260_io_x1 = m_702_io_cout; // @[MUL.scala 253:22]
  assign m_1260_io_x2 = m_709_io_s; // @[MUL.scala 252:21]
  assign m_1260_io_x3 = m_703_io_cout; // @[MUL.scala 253:22]
  assign m_1261_io_x1 = m_710_io_s; // @[MUL.scala 252:21]
  assign m_1261_io_x2 = m_704_io_cout; // @[MUL.scala 253:22]
  assign m_1261_io_x3 = m_711_io_s; // @[MUL.scala 252:21]
  assign m_1262_io_x1 = m_705_io_cout; // @[MUL.scala 253:22]
  assign m_1262_io_x2 = m_712_io_out_0; // @[MUL.scala 104:13]
  assign m_1262_io_x3 = m_706_io_out_1; // @[MUL.scala 105:13]
  assign m_1263_io_x1 = m_713_io_s; // @[MUL.scala 252:21]
  assign m_1263_io_x2 = m_707_io_cout; // @[MUL.scala 253:22]
  assign m_1263_io_x3 = m_714_io_s; // @[MUL.scala 252:21]
  assign m_1264_io_x1 = m_708_io_cout; // @[MUL.scala 253:22]
  assign m_1264_io_x2 = m_715_io_s; // @[MUL.scala 252:21]
  assign m_1264_io_x3 = m_709_io_cout; // @[MUL.scala 253:22]
  assign m_1265_io_x1 = m_716_io_s; // @[MUL.scala 252:21]
  assign m_1265_io_x2 = m_710_io_cout; // @[MUL.scala 253:22]
  assign m_1265_io_x3 = m_717_io_s; // @[MUL.scala 252:21]
  assign m_1266_io_x1 = m_711_io_cout; // @[MUL.scala 253:22]
  assign m_1266_io_x2 = r_2052; // @[MUL.scala 104:13]
  assign m_1266_io_x3 = m_712_io_out_1; // @[MUL.scala 105:13]
  assign m_1267_io_x1 = m_718_io_s; // @[MUL.scala 252:21]
  assign m_1267_io_x2 = m_713_io_cout; // @[MUL.scala 253:22]
  assign m_1267_io_x3 = m_719_io_s; // @[MUL.scala 252:21]
  assign m_1268_io_x1 = m_714_io_cout; // @[MUL.scala 253:22]
  assign m_1268_io_x2 = m_720_io_s; // @[MUL.scala 252:21]
  assign m_1268_io_x3 = m_715_io_cout; // @[MUL.scala 253:22]
  assign m_1269_io_x1 = m_721_io_s; // @[MUL.scala 252:21]
  assign m_1269_io_x2 = m_716_io_cout; // @[MUL.scala 253:22]
  assign m_1269_io_x3 = m_722_io_s; // @[MUL.scala 252:21]
  assign m_1270_io_in_0 = m_717_io_cout; // @[MUL.scala 253:22]
  assign m_1270_io_in_1 = r_2068; // @[MUL.scala 126:16]
  assign m_1271_io_x1 = m_723_io_s; // @[MUL.scala 252:21]
  assign m_1271_io_x2 = m_718_io_cout; // @[MUL.scala 253:22]
  assign m_1271_io_x3 = m_724_io_s; // @[MUL.scala 252:21]
  assign m_1272_io_x1 = m_719_io_cout; // @[MUL.scala 253:22]
  assign m_1272_io_x2 = m_725_io_s; // @[MUL.scala 252:21]
  assign m_1272_io_x3 = m_720_io_cout; // @[MUL.scala 253:22]
  assign m_1273_io_x1 = m_726_io_s; // @[MUL.scala 252:21]
  assign m_1273_io_x2 = m_721_io_cout; // @[MUL.scala 253:22]
  assign m_1273_io_x3 = m_727_io_s; // @[MUL.scala 252:21]
  assign m_1274_io_x1 = m_728_io_s; // @[MUL.scala 252:21]
  assign m_1274_io_x2 = m_723_io_cout; // @[MUL.scala 253:22]
  assign m_1274_io_x3 = m_729_io_s; // @[MUL.scala 252:21]
  assign m_1275_io_x1 = m_724_io_cout; // @[MUL.scala 253:22]
  assign m_1275_io_x2 = m_730_io_s; // @[MUL.scala 252:21]
  assign m_1275_io_x3 = m_725_io_cout; // @[MUL.scala 253:22]
  assign m_1276_io_x1 = m_731_io_s; // @[MUL.scala 252:21]
  assign m_1276_io_x2 = m_726_io_cout; // @[MUL.scala 253:22]
  assign m_1276_io_x3 = m_732_io_s; // @[MUL.scala 252:21]
  assign m_1277_io_x1 = m_733_io_s; // @[MUL.scala 252:21]
  assign m_1277_io_x2 = m_728_io_cout; // @[MUL.scala 253:22]
  assign m_1277_io_x3 = m_734_io_s; // @[MUL.scala 252:21]
  assign m_1278_io_x1 = m_729_io_cout; // @[MUL.scala 253:22]
  assign m_1278_io_x2 = m_735_io_s; // @[MUL.scala 252:21]
  assign m_1278_io_x3 = m_730_io_cout; // @[MUL.scala 253:22]
  assign m_1279_io_x1 = m_736_io_s; // @[MUL.scala 252:21]
  assign m_1279_io_x2 = m_731_io_cout; // @[MUL.scala 253:22]
  assign m_1279_io_x3 = m_737_io_out_0; // @[MUL.scala 105:13]
  assign m_1280_io_x1 = m_738_io_s; // @[MUL.scala 252:21]
  assign m_1280_io_x2 = m_733_io_cout; // @[MUL.scala 253:22]
  assign m_1280_io_x3 = m_739_io_s; // @[MUL.scala 252:21]
  assign m_1281_io_x1 = m_734_io_cout; // @[MUL.scala 253:22]
  assign m_1281_io_x2 = m_740_io_s; // @[MUL.scala 252:21]
  assign m_1281_io_x3 = m_735_io_cout; // @[MUL.scala 253:22]
  assign m_1282_io_x1 = m_741_io_s; // @[MUL.scala 252:21]
  assign m_1282_io_x2 = m_736_io_cout; // @[MUL.scala 253:22]
  assign m_1282_io_x3 = m_742_io_out_0; // @[MUL.scala 105:13]
  assign m_1283_io_x1 = m_743_io_s; // @[MUL.scala 252:21]
  assign m_1283_io_x2 = m_738_io_cout; // @[MUL.scala 253:22]
  assign m_1283_io_x3 = m_744_io_s; // @[MUL.scala 252:21]
  assign m_1284_io_x1 = m_739_io_cout; // @[MUL.scala 253:22]
  assign m_1284_io_x2 = m_745_io_s; // @[MUL.scala 252:21]
  assign m_1284_io_x3 = m_740_io_cout; // @[MUL.scala 253:22]
  assign m_1285_io_x1 = m_746_io_s; // @[MUL.scala 252:21]
  assign m_1285_io_x2 = m_741_io_cout; // @[MUL.scala 253:22]
  assign m_1285_io_x3 = r_2139; // @[MUL.scala 105:13]
  assign m_1286_io_x1 = m_747_io_s; // @[MUL.scala 252:21]
  assign m_1286_io_x2 = m_743_io_cout; // @[MUL.scala 253:22]
  assign m_1286_io_x3 = m_748_io_s; // @[MUL.scala 252:21]
  assign m_1287_io_x1 = m_744_io_cout; // @[MUL.scala 253:22]
  assign m_1287_io_x2 = m_749_io_s; // @[MUL.scala 252:21]
  assign m_1287_io_x3 = m_745_io_cout; // @[MUL.scala 253:22]
  assign m_1288_io_x1 = m_750_io_s; // @[MUL.scala 252:21]
  assign m_1288_io_x2 = m_746_io_cout; // @[MUL.scala 253:22]
  assign m_1288_io_x3 = r_2152; // @[MUL.scala 105:13]
  assign m_1289_io_x1 = m_751_io_s; // @[MUL.scala 252:21]
  assign m_1289_io_x2 = m_747_io_cout; // @[MUL.scala 253:22]
  assign m_1289_io_x3 = m_752_io_s; // @[MUL.scala 252:21]
  assign m_1290_io_x1 = m_748_io_cout; // @[MUL.scala 253:22]
  assign m_1290_io_x2 = m_753_io_s; // @[MUL.scala 252:21]
  assign m_1290_io_x3 = m_749_io_cout; // @[MUL.scala 253:22]
  assign m_1291_io_in_0 = m_754_io_s; // @[MUL.scala 252:21]
  assign m_1291_io_in_1 = m_750_io_cout; // @[MUL.scala 253:22]
  assign m_1292_io_x1 = m_755_io_s; // @[MUL.scala 252:21]
  assign m_1292_io_x2 = m_751_io_cout; // @[MUL.scala 253:22]
  assign m_1292_io_x3 = m_756_io_s; // @[MUL.scala 252:21]
  assign m_1293_io_x1 = m_752_io_cout; // @[MUL.scala 253:22]
  assign m_1293_io_x2 = m_757_io_s; // @[MUL.scala 252:21]
  assign m_1293_io_x3 = m_753_io_cout; // @[MUL.scala 253:22]
  assign m_1294_io_in_0 = m_758_io_s; // @[MUL.scala 252:21]
  assign m_1294_io_in_1 = m_754_io_cout; // @[MUL.scala 253:22]
  assign m_1295_io_x1 = m_759_io_s; // @[MUL.scala 252:21]
  assign m_1295_io_x2 = m_755_io_cout; // @[MUL.scala 253:22]
  assign m_1295_io_x3 = m_760_io_s; // @[MUL.scala 252:21]
  assign m_1296_io_x1 = m_756_io_cout; // @[MUL.scala 253:22]
  assign m_1296_io_x2 = m_761_io_s; // @[MUL.scala 252:21]
  assign m_1296_io_x3 = m_757_io_cout; // @[MUL.scala 253:22]
  assign m_1297_io_in_0 = m_762_io_out_0; // @[MUL.scala 125:16]
  assign m_1297_io_in_1 = m_758_io_cout; // @[MUL.scala 253:22]
  assign m_1298_io_x1 = m_763_io_s; // @[MUL.scala 252:21]
  assign m_1298_io_x2 = m_759_io_cout; // @[MUL.scala 253:22]
  assign m_1298_io_x3 = m_764_io_s; // @[MUL.scala 252:21]
  assign m_1299_io_x1 = m_760_io_cout; // @[MUL.scala 253:22]
  assign m_1299_io_x2 = m_765_io_s; // @[MUL.scala 252:21]
  assign m_1299_io_x3 = m_761_io_cout; // @[MUL.scala 253:22]
  assign m_1300_io_in_0 = m_766_io_out_0; // @[MUL.scala 125:16]
  assign m_1300_io_in_1 = m_762_io_out_1; // @[MUL.scala 126:16]
  assign m_1301_io_x1 = m_767_io_s; // @[MUL.scala 252:21]
  assign m_1301_io_x2 = m_763_io_cout; // @[MUL.scala 253:22]
  assign m_1301_io_x3 = m_768_io_s; // @[MUL.scala 252:21]
  assign m_1302_io_x1 = m_764_io_cout; // @[MUL.scala 253:22]
  assign m_1302_io_x2 = m_769_io_s; // @[MUL.scala 252:21]
  assign m_1302_io_x3 = m_765_io_cout; // @[MUL.scala 253:22]
  assign m_1303_io_in_0 = r_2208; // @[MUL.scala 125:16]
  assign m_1303_io_in_1 = m_766_io_out_1; // @[MUL.scala 126:16]
  assign m_1304_io_x1 = m_770_io_s; // @[MUL.scala 252:21]
  assign m_1304_io_x2 = m_767_io_cout; // @[MUL.scala 253:22]
  assign m_1304_io_x3 = m_771_io_s; // @[MUL.scala 252:21]
  assign m_1305_io_x1 = m_768_io_cout; // @[MUL.scala 253:22]
  assign m_1305_io_x2 = m_772_io_s; // @[MUL.scala 252:21]
  assign m_1305_io_x3 = m_769_io_cout; // @[MUL.scala 253:22]
  assign m_1306_io_x1 = m_773_io_s; // @[MUL.scala 252:21]
  assign m_1306_io_x2 = m_770_io_cout; // @[MUL.scala 253:22]
  assign m_1306_io_x3 = m_774_io_s; // @[MUL.scala 252:21]
  assign m_1307_io_x1 = m_771_io_cout; // @[MUL.scala 253:22]
  assign m_1307_io_x2 = m_775_io_s; // @[MUL.scala 252:21]
  assign m_1307_io_x3 = m_772_io_cout; // @[MUL.scala 253:22]
  assign m_1308_io_x1 = m_776_io_s; // @[MUL.scala 252:21]
  assign m_1308_io_x2 = m_773_io_cout; // @[MUL.scala 253:22]
  assign m_1308_io_x3 = m_777_io_s; // @[MUL.scala 252:21]
  assign m_1309_io_x1 = m_774_io_cout; // @[MUL.scala 253:22]
  assign m_1309_io_x2 = m_778_io_s; // @[MUL.scala 252:21]
  assign m_1309_io_x3 = m_775_io_cout; // @[MUL.scala 253:22]
  assign m_1310_io_x1 = m_779_io_s; // @[MUL.scala 252:21]
  assign m_1310_io_x2 = m_776_io_cout; // @[MUL.scala 253:22]
  assign m_1310_io_x3 = m_780_io_s; // @[MUL.scala 252:21]
  assign m_1311_io_x1 = m_777_io_cout; // @[MUL.scala 253:22]
  assign m_1311_io_x2 = m_781_io_out_0; // @[MUL.scala 104:13]
  assign m_1311_io_x3 = m_778_io_cout; // @[MUL.scala 253:22]
  assign m_1312_io_x1 = m_782_io_s; // @[MUL.scala 252:21]
  assign m_1312_io_x2 = m_779_io_cout; // @[MUL.scala 253:22]
  assign m_1312_io_x3 = m_783_io_s; // @[MUL.scala 252:21]
  assign m_1313_io_x1 = m_780_io_cout; // @[MUL.scala 253:22]
  assign m_1313_io_x2 = m_784_io_out_0; // @[MUL.scala 104:13]
  assign m_1313_io_x3 = m_781_io_out_1; // @[MUL.scala 105:13]
  assign m_1314_io_x1 = m_785_io_s; // @[MUL.scala 252:21]
  assign m_1314_io_x2 = m_782_io_cout; // @[MUL.scala 253:22]
  assign m_1314_io_x3 = m_786_io_s; // @[MUL.scala 252:21]
  assign m_1315_io_x1 = m_783_io_cout; // @[MUL.scala 253:22]
  assign m_1315_io_x2 = r_2259; // @[MUL.scala 104:13]
  assign m_1315_io_x3 = m_784_io_out_1; // @[MUL.scala 105:13]
  assign m_1316_io_x1 = m_787_io_s; // @[MUL.scala 252:21]
  assign m_1316_io_x2 = m_785_io_cout; // @[MUL.scala 253:22]
  assign m_1316_io_x3 = m_788_io_s; // @[MUL.scala 252:21]
  assign m_1317_io_in_0 = m_786_io_cout; // @[MUL.scala 253:22]
  assign m_1317_io_in_1 = r_2266; // @[MUL.scala 126:16]
  assign m_1318_io_x1 = m_789_io_s; // @[MUL.scala 252:21]
  assign m_1318_io_x2 = m_787_io_cout; // @[MUL.scala 253:22]
  assign m_1318_io_x3 = m_790_io_s; // @[MUL.scala 252:21]
  assign m_1319_io_x1 = m_791_io_s; // @[MUL.scala 252:21]
  assign m_1319_io_x2 = m_789_io_cout; // @[MUL.scala 253:22]
  assign m_1319_io_x3 = m_792_io_s; // @[MUL.scala 252:21]
  assign m_1320_io_x1 = m_793_io_s; // @[MUL.scala 252:21]
  assign m_1320_io_x2 = m_791_io_cout; // @[MUL.scala 253:22]
  assign m_1320_io_x3 = m_794_io_out_0; // @[MUL.scala 105:13]
  assign m_1321_io_x1 = m_795_io_s; // @[MUL.scala 252:21]
  assign m_1321_io_x2 = m_793_io_cout; // @[MUL.scala 253:22]
  assign m_1321_io_x3 = m_796_io_out_0; // @[MUL.scala 105:13]
  assign m_1322_io_x1 = m_797_io_s; // @[MUL.scala 252:21]
  assign m_1322_io_x2 = m_795_io_cout; // @[MUL.scala 253:22]
  assign m_1322_io_x3 = r_2292; // @[MUL.scala 105:13]
  assign m_1323_io_x1 = m_798_io_s; // @[MUL.scala 252:21]
  assign m_1323_io_x2 = m_797_io_cout; // @[MUL.scala 253:22]
  assign m_1323_io_x3 = r_2296; // @[MUL.scala 105:13]
  assign m_1324_io_in_0 = m_799_io_s; // @[MUL.scala 252:21]
  assign m_1324_io_in_1 = m_798_io_cout; // @[MUL.scala 253:22]
  assign m_1325_io_in_0 = m_800_io_s; // @[MUL.scala 252:21]
  assign m_1325_io_in_1 = m_799_io_cout; // @[MUL.scala 253:22]
  assign m_1326_io_in_0 = m_801_io_out_0; // @[MUL.scala 125:16]
  assign m_1326_io_in_1 = m_800_io_cout; // @[MUL.scala 253:22]
  assign m_1327_io_in_0 = m_802_io_out_0; // @[MUL.scala 125:16]
  assign m_1327_io_in_1 = m_801_io_out_1; // @[MUL.scala 126:16]
  assign m_1328_io_in_0 = r_2307; // @[MUL.scala 125:16]
  assign m_1328_io_in_1 = m_802_io_out_1; // @[MUL.scala 126:16]
  assign m_1329_io_in_0 = m_804_io_out_0; // @[MUL.scala 125:16]
  assign m_1329_io_in_1 = m_803_io_out_1; // @[MUL.scala 126:16]
  assign m_1330_io_in_0 = m_805_io_out_0; // @[MUL.scala 125:16]
  assign m_1330_io_in_1 = m_804_io_out_1; // @[MUL.scala 126:16]
  assign m_1331_io_in_0 = m_806_io_s; // @[MUL.scala 252:21]
  assign m_1331_io_in_1 = m_805_io_out_1; // @[MUL.scala 126:16]
  assign m_1332_io_in_0 = m_807_io_s; // @[MUL.scala 252:21]
  assign m_1332_io_in_1 = m_806_io_cout; // @[MUL.scala 253:22]
  assign m_1333_io_in_0 = m_808_io_s; // @[MUL.scala 252:21]
  assign m_1333_io_in_1 = m_807_io_cout; // @[MUL.scala 253:22]
  assign m_1334_io_x1 = m_809_io_s; // @[MUL.scala 252:21]
  assign m_1334_io_x2 = m_808_io_cout; // @[MUL.scala 253:22]
  assign m_1334_io_x3 = m_40_io_out_1; // @[MUL.scala 105:13]
  assign m_1335_io_x1 = m_810_io_s; // @[MUL.scala 252:21]
  assign m_1335_io_x2 = m_809_io_cout; // @[MUL.scala 253:22]
  assign m_1335_io_x3 = m_42_io_out_1; // @[MUL.scala 105:13]
  assign m_1336_io_x1 = m_811_io_s; // @[MUL.scala 252:21]
  assign m_1336_io_x2 = m_810_io_cout; // @[MUL.scala 253:22]
  assign m_1336_io_x3 = m_44_io_cout; // @[MUL.scala 253:22]
  assign m_1337_io_x1 = m_812_io_s; // @[MUL.scala 252:21]
  assign m_1337_io_x2 = m_811_io_cout; // @[MUL.scala 253:22]
  assign m_1337_io_x3 = m_813_io_out_0; // @[MUL.scala 105:13]
  assign m_1338_io_x1 = m_814_io_s; // @[MUL.scala 252:21]
  assign m_1338_io_x2 = m_812_io_cout; // @[MUL.scala 253:22]
  assign m_1338_io_x3 = m_815_io_out_0; // @[MUL.scala 105:13]
  assign m_1339_io_x1 = m_816_io_s; // @[MUL.scala 252:21]
  assign m_1339_io_x2 = m_814_io_cout; // @[MUL.scala 253:22]
  assign m_1339_io_x3 = m_817_io_out_0; // @[MUL.scala 105:13]
  assign m_1340_io_x1 = m_818_io_s; // @[MUL.scala 252:21]
  assign m_1340_io_x2 = m_816_io_cout; // @[MUL.scala 253:22]
  assign m_1340_io_x3 = m_819_io_s; // @[MUL.scala 252:21]
  assign m_1341_io_x1 = m_820_io_s; // @[MUL.scala 252:21]
  assign m_1341_io_x2 = m_818_io_cout; // @[MUL.scala 253:22]
  assign m_1341_io_x3 = m_821_io_s; // @[MUL.scala 252:21]
  assign m_1342_io_x1 = m_822_io_s; // @[MUL.scala 252:21]
  assign m_1342_io_x2 = m_820_io_cout; // @[MUL.scala 253:22]
  assign m_1342_io_x3 = m_823_io_s; // @[MUL.scala 252:21]
  assign m_1343_io_x1 = m_824_io_s; // @[MUL.scala 252:21]
  assign m_1343_io_x2 = m_822_io_cout; // @[MUL.scala 253:22]
  assign m_1343_io_x3 = m_825_io_s; // @[MUL.scala 252:21]
  assign m_1344_io_in_0 = m_823_io_cout; // @[MUL.scala 253:22]
  assign m_1344_io_in_1 = r_97; // @[MUL.scala 126:16]
  assign m_1345_io_x1 = m_826_io_s; // @[MUL.scala 252:21]
  assign m_1345_io_x2 = m_824_io_cout; // @[MUL.scala 253:22]
  assign m_1345_io_x3 = m_827_io_s; // @[MUL.scala 252:21]
  assign m_1346_io_in_0 = m_825_io_cout; // @[MUL.scala 253:22]
  assign m_1346_io_in_1 = r_107; // @[MUL.scala 126:16]
  assign m_1347_io_x1 = m_828_io_s; // @[MUL.scala 252:21]
  assign m_1347_io_x2 = m_826_io_cout; // @[MUL.scala 253:22]
  assign m_1347_io_x3 = m_829_io_s; // @[MUL.scala 252:21]
  assign m_1348_io_in_0 = m_827_io_cout; // @[MUL.scala 253:22]
  assign m_1348_io_in_1 = m_72_io_out_0; // @[MUL.scala 126:16]
  assign m_1349_io_x1 = m_830_io_s; // @[MUL.scala 252:21]
  assign m_1349_io_x2 = m_828_io_cout; // @[MUL.scala 253:22]
  assign m_1349_io_x3 = m_831_io_s; // @[MUL.scala 252:21]
  assign m_1350_io_in_0 = m_829_io_cout; // @[MUL.scala 253:22]
  assign m_1350_io_in_1 = m_832_io_out_0; // @[MUL.scala 126:16]
  assign m_1351_io_x1 = m_833_io_s; // @[MUL.scala 252:21]
  assign m_1351_io_x2 = m_830_io_cout; // @[MUL.scala 253:22]
  assign m_1351_io_x3 = m_834_io_s; // @[MUL.scala 252:21]
  assign m_1352_io_x1 = m_831_io_cout; // @[MUL.scala 253:22]
  assign m_1352_io_x2 = m_835_io_out_0; // @[MUL.scala 104:13]
  assign m_1352_io_x3 = m_832_io_out_1; // @[MUL.scala 105:13]
  assign m_1353_io_x1 = m_836_io_s; // @[MUL.scala 252:21]
  assign m_1353_io_x2 = m_833_io_cout; // @[MUL.scala 253:22]
  assign m_1353_io_x3 = m_837_io_s; // @[MUL.scala 252:21]
  assign m_1354_io_x1 = m_834_io_cout; // @[MUL.scala 253:22]
  assign m_1354_io_x2 = m_838_io_out_0; // @[MUL.scala 104:13]
  assign m_1354_io_x3 = m_835_io_out_1; // @[MUL.scala 105:13]
  assign m_1355_io_x1 = m_839_io_s; // @[MUL.scala 252:21]
  assign m_1355_io_x2 = m_836_io_cout; // @[MUL.scala 253:22]
  assign m_1355_io_x3 = m_840_io_s; // @[MUL.scala 252:21]
  assign m_1356_io_x1 = m_837_io_cout; // @[MUL.scala 253:22]
  assign m_1356_io_x2 = m_841_io_s; // @[MUL.scala 252:21]
  assign m_1356_io_x3 = m_838_io_out_1; // @[MUL.scala 105:13]
  assign m_1357_io_x1 = m_842_io_s; // @[MUL.scala 252:21]
  assign m_1357_io_x2 = m_839_io_cout; // @[MUL.scala 253:22]
  assign m_1357_io_x3 = m_843_io_s; // @[MUL.scala 252:21]
  assign m_1358_io_x1 = m_840_io_cout; // @[MUL.scala 253:22]
  assign m_1358_io_x2 = m_844_io_s; // @[MUL.scala 252:21]
  assign m_1358_io_x3 = m_841_io_cout; // @[MUL.scala 253:22]
  assign m_1359_io_x1 = m_845_io_s; // @[MUL.scala 252:21]
  assign m_1359_io_x2 = m_842_io_cout; // @[MUL.scala 253:22]
  assign m_1359_io_x3 = m_846_io_s; // @[MUL.scala 252:21]
  assign m_1360_io_x1 = m_843_io_cout; // @[MUL.scala 253:22]
  assign m_1360_io_x2 = m_847_io_s; // @[MUL.scala 252:21]
  assign m_1360_io_x3 = m_844_io_cout; // @[MUL.scala 253:22]
  assign m_1361_io_x1 = m_848_io_s; // @[MUL.scala 252:21]
  assign m_1361_io_x2 = m_845_io_cout; // @[MUL.scala 253:22]
  assign m_1361_io_x3 = m_849_io_s; // @[MUL.scala 252:21]
  assign m_1362_io_x1 = m_846_io_cout; // @[MUL.scala 253:22]
  assign m_1362_io_x2 = m_850_io_s; // @[MUL.scala 252:21]
  assign m_1362_io_x3 = m_847_io_cout; // @[MUL.scala 253:22]
  assign m_1363_io_x1 = m_851_io_s; // @[MUL.scala 252:21]
  assign m_1363_io_x2 = m_848_io_cout; // @[MUL.scala 253:22]
  assign m_1363_io_x3 = m_852_io_s; // @[MUL.scala 252:21]
  assign m_1364_io_x1 = m_849_io_cout; // @[MUL.scala 253:22]
  assign m_1364_io_x2 = m_853_io_s; // @[MUL.scala 252:21]
  assign m_1364_io_x3 = m_850_io_cout; // @[MUL.scala 253:22]
  assign m_1365_io_x1 = m_854_io_s; // @[MUL.scala 252:21]
  assign m_1365_io_x2 = m_851_io_cout; // @[MUL.scala 253:22]
  assign m_1365_io_x3 = m_855_io_s; // @[MUL.scala 252:21]
  assign m_1366_io_x1 = m_852_io_cout; // @[MUL.scala 253:22]
  assign m_1366_io_x2 = m_856_io_s; // @[MUL.scala 252:21]
  assign m_1366_io_x3 = m_853_io_cout; // @[MUL.scala 253:22]
  assign m_1367_io_x1 = m_857_io_s; // @[MUL.scala 252:21]
  assign m_1367_io_x2 = m_854_io_cout; // @[MUL.scala 253:22]
  assign m_1367_io_x3 = m_858_io_s; // @[MUL.scala 252:21]
  assign m_1368_io_x1 = m_855_io_cout; // @[MUL.scala 253:22]
  assign m_1368_io_x2 = m_859_io_s; // @[MUL.scala 252:21]
  assign m_1368_io_x3 = m_856_io_cout; // @[MUL.scala 253:22]
  assign m_1369_io_x1 = m_861_io_s; // @[MUL.scala 252:21]
  assign m_1369_io_x2 = m_857_io_cout; // @[MUL.scala 253:22]
  assign m_1369_io_x3 = m_862_io_s; // @[MUL.scala 252:21]
  assign m_1370_io_x1 = m_858_io_cout; // @[MUL.scala 253:22]
  assign m_1370_io_x2 = m_863_io_s; // @[MUL.scala 252:21]
  assign m_1370_io_x3 = m_859_io_cout; // @[MUL.scala 253:22]
  assign m_1371_io_in_0 = m_864_io_out_0; // @[MUL.scala 125:16]
  assign m_1371_io_in_1 = m_860_io_out_1; // @[MUL.scala 126:16]
  assign m_1372_io_x1 = m_865_io_s; // @[MUL.scala 252:21]
  assign m_1372_io_x2 = m_861_io_cout; // @[MUL.scala 253:22]
  assign m_1372_io_x3 = m_866_io_s; // @[MUL.scala 252:21]
  assign m_1373_io_x1 = m_862_io_cout; // @[MUL.scala 253:22]
  assign m_1373_io_x2 = m_867_io_s; // @[MUL.scala 252:21]
  assign m_1373_io_x3 = m_863_io_cout; // @[MUL.scala 253:22]
  assign m_1374_io_in_0 = m_868_io_out_0; // @[MUL.scala 125:16]
  assign m_1374_io_in_1 = m_864_io_out_1; // @[MUL.scala 126:16]
  assign m_1375_io_x1 = m_869_io_s; // @[MUL.scala 252:21]
  assign m_1375_io_x2 = m_865_io_cout; // @[MUL.scala 253:22]
  assign m_1375_io_x3 = m_870_io_s; // @[MUL.scala 252:21]
  assign m_1376_io_x1 = m_866_io_cout; // @[MUL.scala 253:22]
  assign m_1376_io_x2 = m_871_io_s; // @[MUL.scala 252:21]
  assign m_1376_io_x3 = m_867_io_cout; // @[MUL.scala 253:22]
  assign m_1377_io_in_0 = m_872_io_s; // @[MUL.scala 252:21]
  assign m_1377_io_in_1 = m_868_io_out_1; // @[MUL.scala 126:16]
  assign m_1378_io_x1 = m_873_io_s; // @[MUL.scala 252:21]
  assign m_1378_io_x2 = m_869_io_cout; // @[MUL.scala 253:22]
  assign m_1378_io_x3 = m_874_io_s; // @[MUL.scala 252:21]
  assign m_1379_io_x1 = m_870_io_cout; // @[MUL.scala 253:22]
  assign m_1379_io_x2 = m_875_io_s; // @[MUL.scala 252:21]
  assign m_1379_io_x3 = m_871_io_cout; // @[MUL.scala 253:22]
  assign m_1380_io_in_0 = m_876_io_s; // @[MUL.scala 252:21]
  assign m_1380_io_in_1 = m_872_io_cout; // @[MUL.scala 253:22]
  assign m_1381_io_x1 = m_877_io_s; // @[MUL.scala 252:21]
  assign m_1381_io_x2 = m_873_io_cout; // @[MUL.scala 253:22]
  assign m_1381_io_x3 = m_878_io_s; // @[MUL.scala 252:21]
  assign m_1382_io_x1 = m_874_io_cout; // @[MUL.scala 253:22]
  assign m_1382_io_x2 = m_879_io_s; // @[MUL.scala 252:21]
  assign m_1382_io_x3 = m_875_io_cout; // @[MUL.scala 253:22]
  assign m_1383_io_in_0 = m_880_io_s; // @[MUL.scala 252:21]
  assign m_1383_io_in_1 = m_876_io_cout; // @[MUL.scala 253:22]
  assign m_1384_io_x1 = m_881_io_s; // @[MUL.scala 252:21]
  assign m_1384_io_x2 = m_877_io_cout; // @[MUL.scala 253:22]
  assign m_1384_io_x3 = m_882_io_s; // @[MUL.scala 252:21]
  assign m_1385_io_x1 = m_878_io_cout; // @[MUL.scala 253:22]
  assign m_1385_io_x2 = m_883_io_s; // @[MUL.scala 252:21]
  assign m_1385_io_x3 = m_879_io_cout; // @[MUL.scala 253:22]
  assign m_1386_io_x1 = m_884_io_s; // @[MUL.scala 252:21]
  assign m_1386_io_x2 = m_880_io_cout; // @[MUL.scala 253:22]
  assign m_1386_io_x3 = r_358; // @[MUL.scala 105:13]
  assign m_1387_io_x1 = m_885_io_s; // @[MUL.scala 252:21]
  assign m_1387_io_x2 = m_881_io_cout; // @[MUL.scala 253:22]
  assign m_1387_io_x3 = m_886_io_s; // @[MUL.scala 252:21]
  assign m_1388_io_x1 = m_882_io_cout; // @[MUL.scala 253:22]
  assign m_1388_io_x2 = m_887_io_s; // @[MUL.scala 252:21]
  assign m_1388_io_x3 = m_883_io_cout; // @[MUL.scala 253:22]
  assign m_1389_io_x1 = m_888_io_s; // @[MUL.scala 252:21]
  assign m_1389_io_x2 = m_884_io_cout; // @[MUL.scala 253:22]
  assign m_1389_io_x3 = r_377; // @[MUL.scala 105:13]
  assign m_1390_io_x1 = m_889_io_s; // @[MUL.scala 252:21]
  assign m_1390_io_x2 = m_885_io_cout; // @[MUL.scala 253:22]
  assign m_1390_io_x3 = m_890_io_s; // @[MUL.scala 252:21]
  assign m_1391_io_x1 = m_886_io_cout; // @[MUL.scala 253:22]
  assign m_1391_io_x2 = m_891_io_s; // @[MUL.scala 252:21]
  assign m_1391_io_x3 = m_887_io_cout; // @[MUL.scala 253:22]
  assign m_1392_io_x1 = m_892_io_s; // @[MUL.scala 252:21]
  assign m_1392_io_x2 = m_888_io_cout; // @[MUL.scala 253:22]
  assign m_1392_io_x3 = m_165_io_out_0; // @[MUL.scala 105:13]
  assign m_1393_io_x1 = m_893_io_s; // @[MUL.scala 252:21]
  assign m_1393_io_x2 = m_889_io_cout; // @[MUL.scala 253:22]
  assign m_1393_io_x3 = m_894_io_s; // @[MUL.scala 252:21]
  assign m_1394_io_x1 = m_890_io_cout; // @[MUL.scala 253:22]
  assign m_1394_io_x2 = m_895_io_s; // @[MUL.scala 252:21]
  assign m_1394_io_x3 = m_891_io_cout; // @[MUL.scala 253:22]
  assign m_1395_io_x1 = m_896_io_s; // @[MUL.scala 252:21]
  assign m_1395_io_x2 = m_892_io_cout; // @[MUL.scala 253:22]
  assign m_1395_io_x3 = m_897_io_out_0; // @[MUL.scala 105:13]
  assign m_1396_io_x1 = m_898_io_s; // @[MUL.scala 252:21]
  assign m_1396_io_x2 = m_893_io_cout; // @[MUL.scala 253:22]
  assign m_1396_io_x3 = m_899_io_s; // @[MUL.scala 252:21]
  assign m_1397_io_x1 = m_894_io_cout; // @[MUL.scala 253:22]
  assign m_1397_io_x2 = m_900_io_s; // @[MUL.scala 252:21]
  assign m_1397_io_x3 = m_895_io_cout; // @[MUL.scala 253:22]
  assign m_1398_io_x1 = m_901_io_s; // @[MUL.scala 252:21]
  assign m_1398_io_x2 = m_896_io_cout; // @[MUL.scala 253:22]
  assign m_1398_io_x3 = m_902_io_out_0; // @[MUL.scala 105:13]
  assign m_1399_io_x1 = m_903_io_s; // @[MUL.scala 252:21]
  assign m_1399_io_x2 = m_898_io_cout; // @[MUL.scala 253:22]
  assign m_1399_io_x3 = m_904_io_s; // @[MUL.scala 252:21]
  assign m_1400_io_x1 = m_899_io_cout; // @[MUL.scala 253:22]
  assign m_1400_io_x2 = m_905_io_s; // @[MUL.scala 252:21]
  assign m_1400_io_x3 = m_900_io_cout; // @[MUL.scala 253:22]
  assign m_1401_io_x1 = m_906_io_s; // @[MUL.scala 252:21]
  assign m_1401_io_x2 = m_901_io_cout; // @[MUL.scala 253:22]
  assign m_1401_io_x3 = m_907_io_out_0; // @[MUL.scala 105:13]
  assign m_1402_io_x1 = m_908_io_s; // @[MUL.scala 252:21]
  assign m_1402_io_x2 = m_903_io_cout; // @[MUL.scala 253:22]
  assign m_1402_io_x3 = m_909_io_s; // @[MUL.scala 252:21]
  assign m_1403_io_x1 = m_904_io_cout; // @[MUL.scala 253:22]
  assign m_1403_io_x2 = m_910_io_s; // @[MUL.scala 252:21]
  assign m_1403_io_x3 = m_905_io_cout; // @[MUL.scala 253:22]
  assign m_1404_io_x1 = m_911_io_s; // @[MUL.scala 252:21]
  assign m_1404_io_x2 = m_906_io_cout; // @[MUL.scala 253:22]
  assign m_1404_io_x3 = m_912_io_s; // @[MUL.scala 252:21]
  assign m_1405_io_x1 = m_913_io_s; // @[MUL.scala 252:21]
  assign m_1405_io_x2 = m_908_io_cout; // @[MUL.scala 253:22]
  assign m_1405_io_x3 = m_914_io_s; // @[MUL.scala 252:21]
  assign m_1406_io_x1 = m_909_io_cout; // @[MUL.scala 253:22]
  assign m_1406_io_x2 = m_915_io_s; // @[MUL.scala 252:21]
  assign m_1406_io_x3 = m_910_io_cout; // @[MUL.scala 253:22]
  assign m_1407_io_x1 = m_916_io_s; // @[MUL.scala 252:21]
  assign m_1407_io_x2 = m_911_io_cout; // @[MUL.scala 253:22]
  assign m_1407_io_x3 = m_917_io_s; // @[MUL.scala 252:21]
  assign m_1408_io_x1 = m_918_io_s; // @[MUL.scala 252:21]
  assign m_1408_io_x2 = m_913_io_cout; // @[MUL.scala 253:22]
  assign m_1408_io_x3 = m_919_io_s; // @[MUL.scala 252:21]
  assign m_1409_io_x1 = m_914_io_cout; // @[MUL.scala 253:22]
  assign m_1409_io_x2 = m_920_io_s; // @[MUL.scala 252:21]
  assign m_1409_io_x3 = m_915_io_cout; // @[MUL.scala 253:22]
  assign m_1410_io_x1 = m_921_io_s; // @[MUL.scala 252:21]
  assign m_1410_io_x2 = m_916_io_cout; // @[MUL.scala 253:22]
  assign m_1410_io_x3 = m_922_io_s; // @[MUL.scala 252:21]
  assign m_1411_io_x1 = m_923_io_s; // @[MUL.scala 252:21]
  assign m_1411_io_x2 = m_918_io_cout; // @[MUL.scala 253:22]
  assign m_1411_io_x3 = m_924_io_s; // @[MUL.scala 252:21]
  assign m_1412_io_x1 = m_919_io_cout; // @[MUL.scala 253:22]
  assign m_1412_io_x2 = m_925_io_s; // @[MUL.scala 252:21]
  assign m_1412_io_x3 = m_920_io_cout; // @[MUL.scala 253:22]
  assign m_1413_io_x1 = m_926_io_s; // @[MUL.scala 252:21]
  assign m_1413_io_x2 = m_921_io_cout; // @[MUL.scala 253:22]
  assign m_1413_io_x3 = m_927_io_s; // @[MUL.scala 252:21]
  assign m_1414_io_in_0 = m_922_io_cout; // @[MUL.scala 253:22]
  assign m_1414_io_in_1 = m_208_io_out_1; // @[MUL.scala 126:16]
  assign m_1415_io_x1 = m_928_io_s; // @[MUL.scala 252:21]
  assign m_1415_io_x2 = m_923_io_cout; // @[MUL.scala 253:22]
  assign m_1415_io_x3 = m_929_io_s; // @[MUL.scala 252:21]
  assign m_1416_io_x1 = m_924_io_cout; // @[MUL.scala 253:22]
  assign m_1416_io_x2 = m_930_io_s; // @[MUL.scala 252:21]
  assign m_1416_io_x3 = m_925_io_cout; // @[MUL.scala 253:22]
  assign m_1417_io_x1 = m_931_io_s; // @[MUL.scala 252:21]
  assign m_1417_io_x2 = m_926_io_cout; // @[MUL.scala 253:22]
  assign m_1417_io_x3 = m_932_io_s; // @[MUL.scala 252:21]
  assign m_1418_io_in_0 = m_927_io_cout; // @[MUL.scala 253:22]
  assign m_1418_io_in_1 = m_216_io_out_1; // @[MUL.scala 126:16]
  assign m_1419_io_x1 = m_933_io_s; // @[MUL.scala 252:21]
  assign m_1419_io_x2 = m_928_io_cout; // @[MUL.scala 253:22]
  assign m_1419_io_x3 = m_934_io_s; // @[MUL.scala 252:21]
  assign m_1420_io_x1 = m_929_io_cout; // @[MUL.scala 253:22]
  assign m_1420_io_x2 = m_935_io_s; // @[MUL.scala 252:21]
  assign m_1420_io_x3 = m_930_io_cout; // @[MUL.scala 253:22]
  assign m_1421_io_x1 = m_936_io_s; // @[MUL.scala 252:21]
  assign m_1421_io_x2 = m_931_io_cout; // @[MUL.scala 253:22]
  assign m_1421_io_x3 = m_937_io_s; // @[MUL.scala 252:21]
  assign m_1422_io_in_0 = m_932_io_cout; // @[MUL.scala 253:22]
  assign m_1422_io_in_1 = m_224_io_cout; // @[MUL.scala 253:22]
  assign m_1423_io_x1 = m_938_io_s; // @[MUL.scala 252:21]
  assign m_1423_io_x2 = m_933_io_cout; // @[MUL.scala 253:22]
  assign m_1423_io_x3 = m_939_io_s; // @[MUL.scala 252:21]
  assign m_1424_io_x1 = m_934_io_cout; // @[MUL.scala 253:22]
  assign m_1424_io_x2 = m_940_io_s; // @[MUL.scala 252:21]
  assign m_1424_io_x3 = m_935_io_cout; // @[MUL.scala 253:22]
  assign m_1425_io_x1 = m_941_io_s; // @[MUL.scala 252:21]
  assign m_1425_io_x2 = m_936_io_cout; // @[MUL.scala 253:22]
  assign m_1425_io_x3 = m_942_io_s; // @[MUL.scala 252:21]
  assign m_1426_io_in_0 = m_937_io_cout; // @[MUL.scala 253:22]
  assign m_1426_io_in_1 = m_943_io_out_0; // @[MUL.scala 126:16]
  assign m_1427_io_x1 = m_944_io_s; // @[MUL.scala 252:21]
  assign m_1427_io_x2 = m_938_io_cout; // @[MUL.scala 253:22]
  assign m_1427_io_x3 = m_945_io_s; // @[MUL.scala 252:21]
  assign m_1428_io_x1 = m_939_io_cout; // @[MUL.scala 253:22]
  assign m_1428_io_x2 = m_946_io_s; // @[MUL.scala 252:21]
  assign m_1428_io_x3 = m_940_io_cout; // @[MUL.scala 253:22]
  assign m_1429_io_x1 = m_947_io_s; // @[MUL.scala 252:21]
  assign m_1429_io_x2 = m_941_io_cout; // @[MUL.scala 253:22]
  assign m_1429_io_x3 = m_948_io_s; // @[MUL.scala 252:21]
  assign m_1430_io_x1 = m_942_io_cout; // @[MUL.scala 253:22]
  assign m_1430_io_x2 = m_949_io_out_0; // @[MUL.scala 104:13]
  assign m_1430_io_x3 = m_943_io_out_1; // @[MUL.scala 105:13]
  assign m_1431_io_x1 = m_950_io_s; // @[MUL.scala 252:21]
  assign m_1431_io_x2 = m_944_io_cout; // @[MUL.scala 253:22]
  assign m_1431_io_x3 = m_951_io_s; // @[MUL.scala 252:21]
  assign m_1432_io_x1 = m_945_io_cout; // @[MUL.scala 253:22]
  assign m_1432_io_x2 = m_952_io_s; // @[MUL.scala 252:21]
  assign m_1432_io_x3 = m_946_io_cout; // @[MUL.scala 253:22]
  assign m_1433_io_x1 = m_953_io_s; // @[MUL.scala 252:21]
  assign m_1433_io_x2 = m_947_io_cout; // @[MUL.scala 253:22]
  assign m_1433_io_x3 = m_954_io_s; // @[MUL.scala 252:21]
  assign m_1434_io_x1 = m_948_io_cout; // @[MUL.scala 253:22]
  assign m_1434_io_x2 = m_955_io_out_0; // @[MUL.scala 104:13]
  assign m_1434_io_x3 = m_949_io_out_1; // @[MUL.scala 105:13]
  assign m_1435_io_x1 = m_956_io_s; // @[MUL.scala 252:21]
  assign m_1435_io_x2 = m_950_io_cout; // @[MUL.scala 253:22]
  assign m_1435_io_x3 = m_957_io_s; // @[MUL.scala 252:21]
  assign m_1436_io_x1 = m_951_io_cout; // @[MUL.scala 253:22]
  assign m_1436_io_x2 = m_958_io_s; // @[MUL.scala 252:21]
  assign m_1436_io_x3 = m_952_io_cout; // @[MUL.scala 253:22]
  assign m_1437_io_x1 = m_959_io_s; // @[MUL.scala 252:21]
  assign m_1437_io_x2 = m_953_io_cout; // @[MUL.scala 253:22]
  assign m_1437_io_x3 = m_960_io_s; // @[MUL.scala 252:21]
  assign m_1438_io_x1 = m_954_io_cout; // @[MUL.scala 253:22]
  assign m_1438_io_x2 = m_961_io_s; // @[MUL.scala 252:21]
  assign m_1438_io_x3 = m_955_io_out_1; // @[MUL.scala 105:13]
  assign m_1439_io_x1 = m_962_io_s; // @[MUL.scala 252:21]
  assign m_1439_io_x2 = m_956_io_cout; // @[MUL.scala 253:22]
  assign m_1439_io_x3 = m_963_io_s; // @[MUL.scala 252:21]
  assign m_1440_io_x1 = m_957_io_cout; // @[MUL.scala 253:22]
  assign m_1440_io_x2 = m_964_io_s; // @[MUL.scala 252:21]
  assign m_1440_io_x3 = m_958_io_cout; // @[MUL.scala 253:22]
  assign m_1441_io_x1 = m_965_io_s; // @[MUL.scala 252:21]
  assign m_1441_io_x2 = m_959_io_cout; // @[MUL.scala 253:22]
  assign m_1441_io_x3 = m_966_io_s; // @[MUL.scala 252:21]
  assign m_1442_io_x1 = m_960_io_cout; // @[MUL.scala 253:22]
  assign m_1442_io_x2 = m_967_io_s; // @[MUL.scala 252:21]
  assign m_1442_io_x3 = m_961_io_cout; // @[MUL.scala 253:22]
  assign m_1443_io_x1 = m_968_io_s; // @[MUL.scala 252:21]
  assign m_1443_io_x2 = m_962_io_cout; // @[MUL.scala 253:22]
  assign m_1443_io_x3 = m_969_io_s; // @[MUL.scala 252:21]
  assign m_1444_io_x1 = m_963_io_cout; // @[MUL.scala 253:22]
  assign m_1444_io_x2 = m_970_io_s; // @[MUL.scala 252:21]
  assign m_1444_io_x3 = m_964_io_cout; // @[MUL.scala 253:22]
  assign m_1445_io_x1 = m_971_io_s; // @[MUL.scala 252:21]
  assign m_1445_io_x2 = m_965_io_cout; // @[MUL.scala 253:22]
  assign m_1445_io_x3 = m_972_io_s; // @[MUL.scala 252:21]
  assign m_1446_io_x1 = m_966_io_cout; // @[MUL.scala 253:22]
  assign m_1446_io_x2 = m_973_io_s; // @[MUL.scala 252:21]
  assign m_1446_io_x3 = m_967_io_cout; // @[MUL.scala 253:22]
  assign m_1447_io_x1 = m_974_io_s; // @[MUL.scala 252:21]
  assign m_1447_io_x2 = m_968_io_cout; // @[MUL.scala 253:22]
  assign m_1447_io_x3 = m_975_io_s; // @[MUL.scala 252:21]
  assign m_1448_io_x1 = m_969_io_cout; // @[MUL.scala 253:22]
  assign m_1448_io_x2 = m_976_io_s; // @[MUL.scala 252:21]
  assign m_1448_io_x3 = m_970_io_cout; // @[MUL.scala 253:22]
  assign m_1449_io_x1 = m_977_io_s; // @[MUL.scala 252:21]
  assign m_1449_io_x2 = m_971_io_cout; // @[MUL.scala 253:22]
  assign m_1449_io_x3 = m_978_io_s; // @[MUL.scala 252:21]
  assign m_1450_io_x1 = m_972_io_cout; // @[MUL.scala 253:22]
  assign m_1450_io_x2 = m_979_io_s; // @[MUL.scala 252:21]
  assign m_1450_io_x3 = m_973_io_cout; // @[MUL.scala 253:22]
  assign m_1451_io_x1 = m_980_io_s; // @[MUL.scala 252:21]
  assign m_1451_io_x2 = m_974_io_cout; // @[MUL.scala 253:22]
  assign m_1451_io_x3 = m_981_io_s; // @[MUL.scala 252:21]
  assign m_1452_io_x1 = m_975_io_cout; // @[MUL.scala 253:22]
  assign m_1452_io_x2 = m_982_io_s; // @[MUL.scala 252:21]
  assign m_1452_io_x3 = m_976_io_cout; // @[MUL.scala 253:22]
  assign m_1453_io_x1 = m_983_io_s; // @[MUL.scala 252:21]
  assign m_1453_io_x2 = m_977_io_cout; // @[MUL.scala 253:22]
  assign m_1453_io_x3 = m_984_io_s; // @[MUL.scala 252:21]
  assign m_1454_io_x1 = m_978_io_cout; // @[MUL.scala 253:22]
  assign m_1454_io_x2 = m_985_io_s; // @[MUL.scala 252:21]
  assign m_1454_io_x3 = m_979_io_cout; // @[MUL.scala 253:22]
  assign m_1455_io_x1 = m_986_io_s; // @[MUL.scala 252:21]
  assign m_1455_io_x2 = m_980_io_cout; // @[MUL.scala 253:22]
  assign m_1455_io_x3 = m_987_io_s; // @[MUL.scala 252:21]
  assign m_1456_io_x1 = m_981_io_cout; // @[MUL.scala 253:22]
  assign m_1456_io_x2 = m_988_io_s; // @[MUL.scala 252:21]
  assign m_1456_io_x3 = m_982_io_cout; // @[MUL.scala 253:22]
  assign m_1457_io_x1 = m_989_io_s; // @[MUL.scala 252:21]
  assign m_1457_io_x2 = m_983_io_cout; // @[MUL.scala 253:22]
  assign m_1457_io_x3 = m_990_io_s; // @[MUL.scala 252:21]
  assign m_1458_io_x1 = m_984_io_cout; // @[MUL.scala 253:22]
  assign m_1458_io_x2 = m_991_io_s; // @[MUL.scala 252:21]
  assign m_1458_io_x3 = m_985_io_cout; // @[MUL.scala 253:22]
  assign m_1459_io_x1 = m_992_io_s; // @[MUL.scala 252:21]
  assign m_1459_io_x2 = m_986_io_cout; // @[MUL.scala 253:22]
  assign m_1459_io_x3 = m_993_io_s; // @[MUL.scala 252:21]
  assign m_1460_io_x1 = m_987_io_cout; // @[MUL.scala 253:22]
  assign m_1460_io_x2 = m_994_io_s; // @[MUL.scala 252:21]
  assign m_1460_io_x3 = m_988_io_cout; // @[MUL.scala 253:22]
  assign m_1461_io_x1 = m_995_io_s; // @[MUL.scala 252:21]
  assign m_1461_io_x2 = m_989_io_cout; // @[MUL.scala 253:22]
  assign m_1461_io_x3 = m_996_io_s; // @[MUL.scala 252:21]
  assign m_1462_io_x1 = m_990_io_cout; // @[MUL.scala 253:22]
  assign m_1462_io_x2 = m_997_io_s; // @[MUL.scala 252:21]
  assign m_1462_io_x3 = m_991_io_cout; // @[MUL.scala 253:22]
  assign m_1463_io_x1 = m_999_io_s; // @[MUL.scala 252:21]
  assign m_1463_io_x2 = m_992_io_cout; // @[MUL.scala 253:22]
  assign m_1463_io_x3 = m_1000_io_s; // @[MUL.scala 252:21]
  assign m_1464_io_x1 = m_993_io_cout; // @[MUL.scala 253:22]
  assign m_1464_io_x2 = m_1001_io_s; // @[MUL.scala 252:21]
  assign m_1464_io_x3 = m_994_io_cout; // @[MUL.scala 253:22]
  assign m_1465_io_x1 = m_1002_io_s; // @[MUL.scala 252:21]
  assign m_1465_io_x2 = m_995_io_cout; // @[MUL.scala 253:22]
  assign m_1465_io_x3 = m_1003_io_s; // @[MUL.scala 252:21]
  assign m_1466_io_x1 = m_996_io_cout; // @[MUL.scala 253:22]
  assign m_1466_io_x2 = m_1004_io_s; // @[MUL.scala 252:21]
  assign m_1466_io_x3 = m_997_io_cout; // @[MUL.scala 253:22]
  assign m_1467_io_in_0 = m_1005_io_out_0; // @[MUL.scala 125:16]
  assign m_1467_io_in_1 = m_998_io_out_1; // @[MUL.scala 126:16]
  assign m_1468_io_x1 = m_1006_io_s; // @[MUL.scala 252:21]
  assign m_1468_io_x2 = m_999_io_cout; // @[MUL.scala 253:22]
  assign m_1468_io_x3 = m_1007_io_s; // @[MUL.scala 252:21]
  assign m_1469_io_x1 = m_1000_io_cout; // @[MUL.scala 253:22]
  assign m_1469_io_x2 = m_1008_io_s; // @[MUL.scala 252:21]
  assign m_1469_io_x3 = m_1001_io_cout; // @[MUL.scala 253:22]
  assign m_1470_io_x1 = m_1009_io_s; // @[MUL.scala 252:21]
  assign m_1470_io_x2 = m_1002_io_cout; // @[MUL.scala 253:22]
  assign m_1470_io_x3 = m_1010_io_s; // @[MUL.scala 252:21]
  assign m_1471_io_x1 = m_1003_io_cout; // @[MUL.scala 253:22]
  assign m_1471_io_x2 = m_1011_io_s; // @[MUL.scala 252:21]
  assign m_1471_io_x3 = m_1004_io_cout; // @[MUL.scala 253:22]
  assign m_1472_io_in_0 = m_1012_io_out_0; // @[MUL.scala 125:16]
  assign m_1472_io_in_1 = m_1005_io_out_1; // @[MUL.scala 126:16]
  assign m_1473_io_x1 = m_1013_io_s; // @[MUL.scala 252:21]
  assign m_1473_io_x2 = m_1006_io_cout; // @[MUL.scala 253:22]
  assign m_1473_io_x3 = m_1014_io_s; // @[MUL.scala 252:21]
  assign m_1474_io_x1 = m_1007_io_cout; // @[MUL.scala 253:22]
  assign m_1474_io_x2 = m_1015_io_s; // @[MUL.scala 252:21]
  assign m_1474_io_x3 = m_1008_io_cout; // @[MUL.scala 253:22]
  assign m_1475_io_x1 = m_1016_io_s; // @[MUL.scala 252:21]
  assign m_1475_io_x2 = m_1009_io_cout; // @[MUL.scala 253:22]
  assign m_1475_io_x3 = m_1017_io_s; // @[MUL.scala 252:21]
  assign m_1476_io_x1 = m_1010_io_cout; // @[MUL.scala 253:22]
  assign m_1476_io_x2 = m_1018_io_s; // @[MUL.scala 252:21]
  assign m_1476_io_x3 = m_1011_io_cout; // @[MUL.scala 253:22]
  assign m_1477_io_in_0 = m_1019_io_s; // @[MUL.scala 252:21]
  assign m_1477_io_in_1 = m_1012_io_out_1; // @[MUL.scala 126:16]
  assign m_1478_io_x1 = m_1020_io_s; // @[MUL.scala 252:21]
  assign m_1478_io_x2 = m_1013_io_cout; // @[MUL.scala 253:22]
  assign m_1478_io_x3 = m_1021_io_s; // @[MUL.scala 252:21]
  assign m_1479_io_x1 = m_1014_io_cout; // @[MUL.scala 253:22]
  assign m_1479_io_x2 = m_1022_io_s; // @[MUL.scala 252:21]
  assign m_1479_io_x3 = m_1015_io_cout; // @[MUL.scala 253:22]
  assign m_1480_io_x1 = m_1023_io_s; // @[MUL.scala 252:21]
  assign m_1480_io_x2 = m_1016_io_cout; // @[MUL.scala 253:22]
  assign m_1480_io_x3 = m_1024_io_s; // @[MUL.scala 252:21]
  assign m_1481_io_x1 = m_1017_io_cout; // @[MUL.scala 253:22]
  assign m_1481_io_x2 = m_1025_io_s; // @[MUL.scala 252:21]
  assign m_1481_io_x3 = m_1018_io_cout; // @[MUL.scala 253:22]
  assign m_1482_io_in_0 = m_1026_io_s; // @[MUL.scala 252:21]
  assign m_1482_io_in_1 = m_1019_io_cout; // @[MUL.scala 253:22]
  assign m_1483_io_x1 = m_1027_io_s; // @[MUL.scala 252:21]
  assign m_1483_io_x2 = m_1020_io_cout; // @[MUL.scala 253:22]
  assign m_1483_io_x3 = m_1028_io_s; // @[MUL.scala 252:21]
  assign m_1484_io_x1 = m_1021_io_cout; // @[MUL.scala 253:22]
  assign m_1484_io_x2 = m_1029_io_s; // @[MUL.scala 252:21]
  assign m_1484_io_x3 = m_1022_io_cout; // @[MUL.scala 253:22]
  assign m_1485_io_x1 = m_1030_io_s; // @[MUL.scala 252:21]
  assign m_1485_io_x2 = m_1023_io_cout; // @[MUL.scala 253:22]
  assign m_1485_io_x3 = m_1031_io_s; // @[MUL.scala 252:21]
  assign m_1486_io_x1 = m_1024_io_cout; // @[MUL.scala 253:22]
  assign m_1486_io_x2 = m_1032_io_s; // @[MUL.scala 252:21]
  assign m_1486_io_x3 = m_1025_io_cout; // @[MUL.scala 253:22]
  assign m_1487_io_in_0 = m_1033_io_s; // @[MUL.scala 252:21]
  assign m_1487_io_in_1 = m_1026_io_cout; // @[MUL.scala 253:22]
  assign m_1488_io_x1 = m_1034_io_s; // @[MUL.scala 252:21]
  assign m_1488_io_x2 = m_1027_io_cout; // @[MUL.scala 253:22]
  assign m_1488_io_x3 = m_1035_io_s; // @[MUL.scala 252:21]
  assign m_1489_io_x1 = m_1028_io_cout; // @[MUL.scala 253:22]
  assign m_1489_io_x2 = m_1036_io_s; // @[MUL.scala 252:21]
  assign m_1489_io_x3 = m_1029_io_cout; // @[MUL.scala 253:22]
  assign m_1490_io_x1 = m_1037_io_s; // @[MUL.scala 252:21]
  assign m_1490_io_x2 = m_1030_io_cout; // @[MUL.scala 253:22]
  assign m_1490_io_x3 = m_1038_io_s; // @[MUL.scala 252:21]
  assign m_1491_io_x1 = m_1031_io_cout; // @[MUL.scala 253:22]
  assign m_1491_io_x2 = m_1039_io_s; // @[MUL.scala 252:21]
  assign m_1491_io_x3 = m_1032_io_cout; // @[MUL.scala 253:22]
  assign m_1492_io_x1 = m_1040_io_s; // @[MUL.scala 252:21]
  assign m_1492_io_x2 = m_1033_io_cout; // @[MUL.scala 253:22]
  assign m_1492_io_x3 = m_373_io_out_1; // @[MUL.scala 105:13]
  assign m_1493_io_x1 = m_1041_io_s; // @[MUL.scala 252:21]
  assign m_1493_io_x2 = m_1034_io_cout; // @[MUL.scala 253:22]
  assign m_1493_io_x3 = m_1042_io_s; // @[MUL.scala 252:21]
  assign m_1494_io_x1 = m_1035_io_cout; // @[MUL.scala 253:22]
  assign m_1494_io_x2 = m_1043_io_s; // @[MUL.scala 252:21]
  assign m_1494_io_x3 = m_1036_io_cout; // @[MUL.scala 253:22]
  assign m_1495_io_x1 = m_1044_io_s; // @[MUL.scala 252:21]
  assign m_1495_io_x2 = m_1037_io_cout; // @[MUL.scala 253:22]
  assign m_1495_io_x3 = m_1045_io_s; // @[MUL.scala 252:21]
  assign m_1496_io_x1 = m_1038_io_cout; // @[MUL.scala 253:22]
  assign m_1496_io_x2 = m_1046_io_s; // @[MUL.scala 252:21]
  assign m_1496_io_x3 = m_1039_io_cout; // @[MUL.scala 253:22]
  assign m_1497_io_x1 = m_1047_io_s; // @[MUL.scala 252:21]
  assign m_1497_io_x2 = m_1040_io_cout; // @[MUL.scala 253:22]
  assign m_1497_io_x3 = m_384_io_out_1; // @[MUL.scala 105:13]
  assign m_1498_io_x1 = m_1048_io_s; // @[MUL.scala 252:21]
  assign m_1498_io_x2 = m_1041_io_cout; // @[MUL.scala 253:22]
  assign m_1498_io_x3 = m_1049_io_s; // @[MUL.scala 252:21]
  assign m_1499_io_x1 = m_1042_io_cout; // @[MUL.scala 253:22]
  assign m_1499_io_x2 = m_1050_io_s; // @[MUL.scala 252:21]
  assign m_1499_io_x3 = m_1043_io_cout; // @[MUL.scala 253:22]
  assign m_1500_io_x1 = m_1051_io_s; // @[MUL.scala 252:21]
  assign m_1500_io_x2 = m_1044_io_cout; // @[MUL.scala 253:22]
  assign m_1500_io_x3 = m_1052_io_s; // @[MUL.scala 252:21]
  assign m_1501_io_x1 = m_1045_io_cout; // @[MUL.scala 253:22]
  assign m_1501_io_x2 = m_1053_io_s; // @[MUL.scala 252:21]
  assign m_1501_io_x3 = m_1046_io_cout; // @[MUL.scala 253:22]
  assign m_1502_io_x1 = m_1054_io_s; // @[MUL.scala 252:21]
  assign m_1502_io_x2 = m_1047_io_cout; // @[MUL.scala 253:22]
  assign m_1502_io_x3 = m_395_io_cout; // @[MUL.scala 253:22]
  assign m_1503_io_x1 = m_1055_io_s; // @[MUL.scala 252:21]
  assign m_1503_io_x2 = m_1048_io_cout; // @[MUL.scala 253:22]
  assign m_1503_io_x3 = m_1056_io_s; // @[MUL.scala 252:21]
  assign m_1504_io_x1 = m_1049_io_cout; // @[MUL.scala 253:22]
  assign m_1504_io_x2 = m_1057_io_s; // @[MUL.scala 252:21]
  assign m_1504_io_x3 = m_1050_io_cout; // @[MUL.scala 253:22]
  assign m_1505_io_x1 = m_1058_io_s; // @[MUL.scala 252:21]
  assign m_1505_io_x2 = m_1051_io_cout; // @[MUL.scala 253:22]
  assign m_1505_io_x3 = m_1059_io_s; // @[MUL.scala 252:21]
  assign m_1506_io_x1 = m_1052_io_cout; // @[MUL.scala 253:22]
  assign m_1506_io_x2 = m_1060_io_s; // @[MUL.scala 252:21]
  assign m_1506_io_x3 = m_1053_io_cout; // @[MUL.scala 253:22]
  assign m_1507_io_x1 = m_1061_io_s; // @[MUL.scala 252:21]
  assign m_1507_io_x2 = m_1054_io_cout; // @[MUL.scala 253:22]
  assign m_1507_io_x3 = m_406_io_cout; // @[MUL.scala 253:22]
  assign m_1508_io_x1 = m_1062_io_s; // @[MUL.scala 252:21]
  assign m_1508_io_x2 = m_1055_io_cout; // @[MUL.scala 253:22]
  assign m_1508_io_x3 = m_1063_io_s; // @[MUL.scala 252:21]
  assign m_1509_io_x1 = m_1056_io_cout; // @[MUL.scala 253:22]
  assign m_1509_io_x2 = m_1064_io_s; // @[MUL.scala 252:21]
  assign m_1509_io_x3 = m_1057_io_cout; // @[MUL.scala 253:22]
  assign m_1510_io_x1 = m_1065_io_s; // @[MUL.scala 252:21]
  assign m_1510_io_x2 = m_1058_io_cout; // @[MUL.scala 253:22]
  assign m_1510_io_x3 = m_1066_io_s; // @[MUL.scala 252:21]
  assign m_1511_io_x1 = m_1059_io_cout; // @[MUL.scala 253:22]
  assign m_1511_io_x2 = m_1067_io_s; // @[MUL.scala 252:21]
  assign m_1511_io_x3 = m_1060_io_cout; // @[MUL.scala 253:22]
  assign m_1512_io_x1 = m_1068_io_s; // @[MUL.scala 252:21]
  assign m_1512_io_x2 = m_1061_io_cout; // @[MUL.scala 253:22]
  assign m_1512_io_x3 = m_417_io_cout; // @[MUL.scala 253:22]
  assign m_1513_io_x1 = m_1069_io_s; // @[MUL.scala 252:21]
  assign m_1513_io_x2 = m_1062_io_cout; // @[MUL.scala 253:22]
  assign m_1513_io_x3 = m_1070_io_s; // @[MUL.scala 252:21]
  assign m_1514_io_x1 = m_1063_io_cout; // @[MUL.scala 253:22]
  assign m_1514_io_x2 = m_1071_io_s; // @[MUL.scala 252:21]
  assign m_1514_io_x3 = m_1064_io_cout; // @[MUL.scala 253:22]
  assign m_1515_io_x1 = m_1072_io_s; // @[MUL.scala 252:21]
  assign m_1515_io_x2 = m_1065_io_cout; // @[MUL.scala 253:22]
  assign m_1515_io_x3 = m_1073_io_s; // @[MUL.scala 252:21]
  assign m_1516_io_x1 = m_1066_io_cout; // @[MUL.scala 253:22]
  assign m_1516_io_x2 = m_1074_io_s; // @[MUL.scala 252:21]
  assign m_1516_io_x3 = m_1067_io_cout; // @[MUL.scala 253:22]
  assign m_1517_io_x1 = m_1075_io_s; // @[MUL.scala 252:21]
  assign m_1517_io_x2 = m_1068_io_cout; // @[MUL.scala 253:22]
  assign m_1517_io_x3 = m_428_io_cout; // @[MUL.scala 253:22]
  assign m_1518_io_x1 = m_1076_io_s; // @[MUL.scala 252:21]
  assign m_1518_io_x2 = m_1069_io_cout; // @[MUL.scala 253:22]
  assign m_1518_io_x3 = m_1077_io_s; // @[MUL.scala 252:21]
  assign m_1519_io_x1 = m_1070_io_cout; // @[MUL.scala 253:22]
  assign m_1519_io_x2 = m_1078_io_s; // @[MUL.scala 252:21]
  assign m_1519_io_x3 = m_1071_io_cout; // @[MUL.scala 253:22]
  assign m_1520_io_x1 = m_1079_io_s; // @[MUL.scala 252:21]
  assign m_1520_io_x2 = m_1072_io_cout; // @[MUL.scala 253:22]
  assign m_1520_io_x3 = m_1080_io_s; // @[MUL.scala 252:21]
  assign m_1521_io_x1 = m_1073_io_cout; // @[MUL.scala 253:22]
  assign m_1521_io_x2 = m_1081_io_s; // @[MUL.scala 252:21]
  assign m_1521_io_x3 = m_1074_io_cout; // @[MUL.scala 253:22]
  assign m_1522_io_x1 = m_1082_io_s; // @[MUL.scala 252:21]
  assign m_1522_io_x2 = m_1075_io_cout; // @[MUL.scala 253:22]
  assign m_1522_io_x3 = m_439_io_cout; // @[MUL.scala 253:22]
  assign m_1523_io_x1 = m_1083_io_s; // @[MUL.scala 252:21]
  assign m_1523_io_x2 = m_1076_io_cout; // @[MUL.scala 253:22]
  assign m_1523_io_x3 = m_1084_io_s; // @[MUL.scala 252:21]
  assign m_1524_io_x1 = m_1077_io_cout; // @[MUL.scala 253:22]
  assign m_1524_io_x2 = m_1085_io_s; // @[MUL.scala 252:21]
  assign m_1524_io_x3 = m_1078_io_cout; // @[MUL.scala 253:22]
  assign m_1525_io_x1 = m_1086_io_s; // @[MUL.scala 252:21]
  assign m_1525_io_x2 = m_1079_io_cout; // @[MUL.scala 253:22]
  assign m_1525_io_x3 = m_1087_io_s; // @[MUL.scala 252:21]
  assign m_1526_io_x1 = m_1080_io_cout; // @[MUL.scala 253:22]
  assign m_1526_io_x2 = m_1088_io_s; // @[MUL.scala 252:21]
  assign m_1526_io_x3 = m_1081_io_cout; // @[MUL.scala 253:22]
  assign m_1527_io_x1 = m_1089_io_s; // @[MUL.scala 252:21]
  assign m_1527_io_x2 = m_1082_io_cout; // @[MUL.scala 253:22]
  assign m_1527_io_x3 = m_450_io_cout; // @[MUL.scala 253:22]
  assign m_1528_io_x1 = m_1090_io_s; // @[MUL.scala 252:21]
  assign m_1528_io_x2 = m_1083_io_cout; // @[MUL.scala 253:22]
  assign m_1528_io_x3 = m_1091_io_s; // @[MUL.scala 252:21]
  assign m_1529_io_x1 = m_1084_io_cout; // @[MUL.scala 253:22]
  assign m_1529_io_x2 = m_1092_io_s; // @[MUL.scala 252:21]
  assign m_1529_io_x3 = m_1085_io_cout; // @[MUL.scala 253:22]
  assign m_1530_io_x1 = m_1093_io_s; // @[MUL.scala 252:21]
  assign m_1530_io_x2 = m_1086_io_cout; // @[MUL.scala 253:22]
  assign m_1530_io_x3 = m_1094_io_s; // @[MUL.scala 252:21]
  assign m_1531_io_x1 = m_1087_io_cout; // @[MUL.scala 253:22]
  assign m_1531_io_x2 = m_1095_io_s; // @[MUL.scala 252:21]
  assign m_1531_io_x3 = m_1088_io_cout; // @[MUL.scala 253:22]
  assign m_1532_io_x1 = m_1096_io_s; // @[MUL.scala 252:21]
  assign m_1532_io_x2 = m_1089_io_cout; // @[MUL.scala 253:22]
  assign m_1532_io_x3 = m_461_io_cout; // @[MUL.scala 253:22]
  assign m_1533_io_x1 = m_1097_io_s; // @[MUL.scala 252:21]
  assign m_1533_io_x2 = m_1090_io_cout; // @[MUL.scala 253:22]
  assign m_1533_io_x3 = m_1098_io_s; // @[MUL.scala 252:21]
  assign m_1534_io_x1 = m_1091_io_cout; // @[MUL.scala 253:22]
  assign m_1534_io_x2 = m_1099_io_s; // @[MUL.scala 252:21]
  assign m_1534_io_x3 = m_1092_io_cout; // @[MUL.scala 253:22]
  assign m_1535_io_x1 = m_1100_io_s; // @[MUL.scala 252:21]
  assign m_1535_io_x2 = m_1093_io_cout; // @[MUL.scala 253:22]
  assign m_1535_io_x3 = m_1101_io_s; // @[MUL.scala 252:21]
  assign m_1536_io_x1 = m_1094_io_cout; // @[MUL.scala 253:22]
  assign m_1536_io_x2 = m_1102_io_s; // @[MUL.scala 252:21]
  assign m_1536_io_x3 = m_1095_io_cout; // @[MUL.scala 253:22]
  assign m_1537_io_x1 = m_1103_io_s; // @[MUL.scala 252:21]
  assign m_1537_io_x2 = m_1096_io_cout; // @[MUL.scala 253:22]
  assign m_1537_io_x3 = m_472_io_out_1; // @[MUL.scala 105:13]
  assign m_1538_io_x1 = m_1104_io_s; // @[MUL.scala 252:21]
  assign m_1538_io_x2 = m_1097_io_cout; // @[MUL.scala 253:22]
  assign m_1538_io_x3 = m_1105_io_s; // @[MUL.scala 252:21]
  assign m_1539_io_x1 = m_1098_io_cout; // @[MUL.scala 253:22]
  assign m_1539_io_x2 = m_1106_io_s; // @[MUL.scala 252:21]
  assign m_1539_io_x3 = m_1099_io_cout; // @[MUL.scala 253:22]
  assign m_1540_io_x1 = m_1107_io_s; // @[MUL.scala 252:21]
  assign m_1540_io_x2 = m_1100_io_cout; // @[MUL.scala 253:22]
  assign m_1540_io_x3 = m_1108_io_s; // @[MUL.scala 252:21]
  assign m_1541_io_x1 = m_1101_io_cout; // @[MUL.scala 253:22]
  assign m_1541_io_x2 = m_1109_io_s; // @[MUL.scala 252:21]
  assign m_1541_io_x3 = m_1102_io_cout; // @[MUL.scala 253:22]
  assign m_1542_io_in_0 = m_1110_io_s; // @[MUL.scala 252:21]
  assign m_1542_io_in_1 = m_1103_io_cout; // @[MUL.scala 253:22]
  assign m_1543_io_x1 = m_1111_io_s; // @[MUL.scala 252:21]
  assign m_1543_io_x2 = m_1104_io_cout; // @[MUL.scala 253:22]
  assign m_1543_io_x3 = m_1112_io_s; // @[MUL.scala 252:21]
  assign m_1544_io_x1 = m_1105_io_cout; // @[MUL.scala 253:22]
  assign m_1544_io_x2 = m_1113_io_s; // @[MUL.scala 252:21]
  assign m_1544_io_x3 = m_1106_io_cout; // @[MUL.scala 253:22]
  assign m_1545_io_x1 = m_1114_io_s; // @[MUL.scala 252:21]
  assign m_1545_io_x2 = m_1107_io_cout; // @[MUL.scala 253:22]
  assign m_1545_io_x3 = m_1115_io_s; // @[MUL.scala 252:21]
  assign m_1546_io_x1 = m_1108_io_cout; // @[MUL.scala 253:22]
  assign m_1546_io_x2 = m_1116_io_s; // @[MUL.scala 252:21]
  assign m_1546_io_x3 = m_1109_io_cout; // @[MUL.scala 253:22]
  assign m_1547_io_in_0 = m_1117_io_out_0; // @[MUL.scala 125:16]
  assign m_1547_io_in_1 = m_1110_io_cout; // @[MUL.scala 253:22]
  assign m_1548_io_x1 = m_1118_io_s; // @[MUL.scala 252:21]
  assign m_1548_io_x2 = m_1111_io_cout; // @[MUL.scala 253:22]
  assign m_1548_io_x3 = m_1119_io_s; // @[MUL.scala 252:21]
  assign m_1549_io_x1 = m_1112_io_cout; // @[MUL.scala 253:22]
  assign m_1549_io_x2 = m_1120_io_s; // @[MUL.scala 252:21]
  assign m_1549_io_x3 = m_1113_io_cout; // @[MUL.scala 253:22]
  assign m_1550_io_x1 = m_1121_io_s; // @[MUL.scala 252:21]
  assign m_1550_io_x2 = m_1114_io_cout; // @[MUL.scala 253:22]
  assign m_1550_io_x3 = m_1122_io_s; // @[MUL.scala 252:21]
  assign m_1551_io_x1 = m_1115_io_cout; // @[MUL.scala 253:22]
  assign m_1551_io_x2 = m_1123_io_s; // @[MUL.scala 252:21]
  assign m_1551_io_x3 = m_1116_io_cout; // @[MUL.scala 253:22]
  assign m_1552_io_in_0 = m_1124_io_out_0; // @[MUL.scala 125:16]
  assign m_1552_io_in_1 = m_1117_io_out_1; // @[MUL.scala 126:16]
  assign m_1553_io_x1 = m_1125_io_s; // @[MUL.scala 252:21]
  assign m_1553_io_x2 = m_1118_io_cout; // @[MUL.scala 253:22]
  assign m_1553_io_x3 = m_1126_io_s; // @[MUL.scala 252:21]
  assign m_1554_io_x1 = m_1119_io_cout; // @[MUL.scala 253:22]
  assign m_1554_io_x2 = m_1127_io_s; // @[MUL.scala 252:21]
  assign m_1554_io_x3 = m_1120_io_cout; // @[MUL.scala 253:22]
  assign m_1555_io_x1 = m_1128_io_s; // @[MUL.scala 252:21]
  assign m_1555_io_x2 = m_1121_io_cout; // @[MUL.scala 253:22]
  assign m_1555_io_x3 = m_1129_io_s; // @[MUL.scala 252:21]
  assign m_1556_io_x1 = m_1122_io_cout; // @[MUL.scala 253:22]
  assign m_1556_io_x2 = m_1130_io_s; // @[MUL.scala 252:21]
  assign m_1556_io_x3 = m_1123_io_cout; // @[MUL.scala 253:22]
  assign m_1557_io_in_0 = m_1131_io_out_0; // @[MUL.scala 125:16]
  assign m_1557_io_in_1 = m_1124_io_out_1; // @[MUL.scala 126:16]
  assign m_1558_io_x1 = m_1132_io_s; // @[MUL.scala 252:21]
  assign m_1558_io_x2 = m_1125_io_cout; // @[MUL.scala 253:22]
  assign m_1558_io_x3 = m_1133_io_s; // @[MUL.scala 252:21]
  assign m_1559_io_x1 = m_1126_io_cout; // @[MUL.scala 253:22]
  assign m_1559_io_x2 = m_1134_io_s; // @[MUL.scala 252:21]
  assign m_1559_io_x3 = m_1127_io_cout; // @[MUL.scala 253:22]
  assign m_1560_io_x1 = m_1135_io_s; // @[MUL.scala 252:21]
  assign m_1560_io_x2 = m_1128_io_cout; // @[MUL.scala 253:22]
  assign m_1560_io_x3 = m_1136_io_s; // @[MUL.scala 252:21]
  assign m_1561_io_x1 = m_1129_io_cout; // @[MUL.scala 253:22]
  assign m_1561_io_x2 = m_1137_io_s; // @[MUL.scala 252:21]
  assign m_1561_io_x3 = m_1130_io_cout; // @[MUL.scala 253:22]
  assign m_1562_io_in_0 = m_1138_io_out_0; // @[MUL.scala 125:16]
  assign m_1562_io_in_1 = m_1131_io_out_1; // @[MUL.scala 126:16]
  assign m_1563_io_x1 = m_1139_io_s; // @[MUL.scala 252:21]
  assign m_1563_io_x2 = m_1132_io_cout; // @[MUL.scala 253:22]
  assign m_1563_io_x3 = m_1140_io_s; // @[MUL.scala 252:21]
  assign m_1564_io_x1 = m_1133_io_cout; // @[MUL.scala 253:22]
  assign m_1564_io_x2 = m_1141_io_s; // @[MUL.scala 252:21]
  assign m_1564_io_x3 = m_1134_io_cout; // @[MUL.scala 253:22]
  assign m_1565_io_x1 = m_1142_io_s; // @[MUL.scala 252:21]
  assign m_1565_io_x2 = m_1135_io_cout; // @[MUL.scala 253:22]
  assign m_1565_io_x3 = m_1143_io_s; // @[MUL.scala 252:21]
  assign m_1566_io_x1 = m_1136_io_cout; // @[MUL.scala 253:22]
  assign m_1566_io_x2 = m_1144_io_s; // @[MUL.scala 252:21]
  assign m_1566_io_x3 = m_1137_io_cout; // @[MUL.scala 253:22]
  assign m_1567_io_in_0 = m_1145_io_out_0; // @[MUL.scala 125:16]
  assign m_1567_io_in_1 = m_1138_io_out_1; // @[MUL.scala 126:16]
  assign m_1568_io_x1 = m_1146_io_s; // @[MUL.scala 252:21]
  assign m_1568_io_x2 = m_1139_io_cout; // @[MUL.scala 253:22]
  assign m_1568_io_x3 = m_1147_io_s; // @[MUL.scala 252:21]
  assign m_1569_io_x1 = m_1140_io_cout; // @[MUL.scala 253:22]
  assign m_1569_io_x2 = m_1148_io_s; // @[MUL.scala 252:21]
  assign m_1569_io_x3 = m_1141_io_cout; // @[MUL.scala 253:22]
  assign m_1570_io_x1 = m_1149_io_s; // @[MUL.scala 252:21]
  assign m_1570_io_x2 = m_1142_io_cout; // @[MUL.scala 253:22]
  assign m_1570_io_x3 = m_1150_io_s; // @[MUL.scala 252:21]
  assign m_1571_io_x1 = m_1143_io_cout; // @[MUL.scala 253:22]
  assign m_1571_io_x2 = m_1151_io_s; // @[MUL.scala 252:21]
  assign m_1571_io_x3 = m_1144_io_cout; // @[MUL.scala 253:22]
  assign m_1572_io_in_0 = r_1552; // @[MUL.scala 125:16]
  assign m_1572_io_in_1 = m_1145_io_out_1; // @[MUL.scala 126:16]
  assign m_1573_io_x1 = m_1152_io_s; // @[MUL.scala 252:21]
  assign m_1573_io_x2 = m_1146_io_cout; // @[MUL.scala 253:22]
  assign m_1573_io_x3 = m_1153_io_s; // @[MUL.scala 252:21]
  assign m_1574_io_x1 = m_1147_io_cout; // @[MUL.scala 253:22]
  assign m_1574_io_x2 = m_1154_io_s; // @[MUL.scala 252:21]
  assign m_1574_io_x3 = m_1148_io_cout; // @[MUL.scala 253:22]
  assign m_1575_io_x1 = m_1155_io_s; // @[MUL.scala 252:21]
  assign m_1575_io_x2 = m_1149_io_cout; // @[MUL.scala 253:22]
  assign m_1575_io_x3 = m_1156_io_s; // @[MUL.scala 252:21]
  assign m_1576_io_x1 = m_1150_io_cout; // @[MUL.scala 253:22]
  assign m_1576_io_x2 = m_1157_io_s; // @[MUL.scala 252:21]
  assign m_1576_io_x3 = m_1151_io_cout; // @[MUL.scala 253:22]
  assign m_1577_io_x1 = m_1158_io_s; // @[MUL.scala 252:21]
  assign m_1577_io_x2 = m_1152_io_cout; // @[MUL.scala 253:22]
  assign m_1577_io_x3 = m_1159_io_s; // @[MUL.scala 252:21]
  assign m_1578_io_x1 = m_1153_io_cout; // @[MUL.scala 253:22]
  assign m_1578_io_x2 = m_1160_io_s; // @[MUL.scala 252:21]
  assign m_1578_io_x3 = m_1154_io_cout; // @[MUL.scala 253:22]
  assign m_1579_io_x1 = m_1161_io_s; // @[MUL.scala 252:21]
  assign m_1579_io_x2 = m_1155_io_cout; // @[MUL.scala 253:22]
  assign m_1579_io_x3 = m_1162_io_s; // @[MUL.scala 252:21]
  assign m_1580_io_x1 = m_1156_io_cout; // @[MUL.scala 253:22]
  assign m_1580_io_x2 = m_1163_io_s; // @[MUL.scala 252:21]
  assign m_1580_io_x3 = m_1157_io_cout; // @[MUL.scala 253:22]
  assign m_1581_io_x1 = m_1164_io_s; // @[MUL.scala 252:21]
  assign m_1581_io_x2 = m_1158_io_cout; // @[MUL.scala 253:22]
  assign m_1581_io_x3 = m_1165_io_s; // @[MUL.scala 252:21]
  assign m_1582_io_x1 = m_1159_io_cout; // @[MUL.scala 253:22]
  assign m_1582_io_x2 = m_1166_io_s; // @[MUL.scala 252:21]
  assign m_1582_io_x3 = m_1160_io_cout; // @[MUL.scala 253:22]
  assign m_1583_io_x1 = m_1167_io_s; // @[MUL.scala 252:21]
  assign m_1583_io_x2 = m_1161_io_cout; // @[MUL.scala 253:22]
  assign m_1583_io_x3 = m_1168_io_s; // @[MUL.scala 252:21]
  assign m_1584_io_x1 = m_1162_io_cout; // @[MUL.scala 253:22]
  assign m_1584_io_x2 = m_1169_io_s; // @[MUL.scala 252:21]
  assign m_1584_io_x3 = m_1163_io_cout; // @[MUL.scala 253:22]
  assign m_1585_io_x1 = m_1170_io_s; // @[MUL.scala 252:21]
  assign m_1585_io_x2 = m_1164_io_cout; // @[MUL.scala 253:22]
  assign m_1585_io_x3 = m_1171_io_s; // @[MUL.scala 252:21]
  assign m_1586_io_x1 = m_1165_io_cout; // @[MUL.scala 253:22]
  assign m_1586_io_x2 = m_1172_io_s; // @[MUL.scala 252:21]
  assign m_1586_io_x3 = m_1166_io_cout; // @[MUL.scala 253:22]
  assign m_1587_io_x1 = m_1173_io_s; // @[MUL.scala 252:21]
  assign m_1587_io_x2 = m_1167_io_cout; // @[MUL.scala 253:22]
  assign m_1587_io_x3 = m_1174_io_s; // @[MUL.scala 252:21]
  assign m_1588_io_x1 = m_1168_io_cout; // @[MUL.scala 253:22]
  assign m_1588_io_x2 = m_1175_io_s; // @[MUL.scala 252:21]
  assign m_1588_io_x3 = m_1169_io_cout; // @[MUL.scala 253:22]
  assign m_1589_io_x1 = m_1176_io_s; // @[MUL.scala 252:21]
  assign m_1589_io_x2 = m_1170_io_cout; // @[MUL.scala 253:22]
  assign m_1589_io_x3 = m_1177_io_s; // @[MUL.scala 252:21]
  assign m_1590_io_x1 = m_1171_io_cout; // @[MUL.scala 253:22]
  assign m_1590_io_x2 = m_1178_io_s; // @[MUL.scala 252:21]
  assign m_1590_io_x3 = m_1172_io_cout; // @[MUL.scala 253:22]
  assign m_1591_io_x1 = m_1179_io_s; // @[MUL.scala 252:21]
  assign m_1591_io_x2 = m_1173_io_cout; // @[MUL.scala 253:22]
  assign m_1591_io_x3 = m_1180_io_s; // @[MUL.scala 252:21]
  assign m_1592_io_x1 = m_1174_io_cout; // @[MUL.scala 253:22]
  assign m_1592_io_x2 = m_1181_io_s; // @[MUL.scala 252:21]
  assign m_1592_io_x3 = m_1175_io_cout; // @[MUL.scala 253:22]
  assign m_1593_io_x1 = m_1182_io_s; // @[MUL.scala 252:21]
  assign m_1593_io_x2 = m_1176_io_cout; // @[MUL.scala 253:22]
  assign m_1593_io_x3 = m_1183_io_s; // @[MUL.scala 252:21]
  assign m_1594_io_x1 = m_1177_io_cout; // @[MUL.scala 253:22]
  assign m_1594_io_x2 = m_1184_io_s; // @[MUL.scala 252:21]
  assign m_1594_io_x3 = m_1178_io_cout; // @[MUL.scala 253:22]
  assign m_1595_io_x1 = m_1185_io_s; // @[MUL.scala 252:21]
  assign m_1595_io_x2 = m_1179_io_cout; // @[MUL.scala 253:22]
  assign m_1595_io_x3 = m_1186_io_s; // @[MUL.scala 252:21]
  assign m_1596_io_x1 = m_1180_io_cout; // @[MUL.scala 253:22]
  assign m_1596_io_x2 = m_1187_io_out_0; // @[MUL.scala 104:13]
  assign m_1596_io_x3 = m_1181_io_cout; // @[MUL.scala 253:22]
  assign m_1597_io_x1 = m_1188_io_s; // @[MUL.scala 252:21]
  assign m_1597_io_x2 = m_1182_io_cout; // @[MUL.scala 253:22]
  assign m_1597_io_x3 = m_1189_io_s; // @[MUL.scala 252:21]
  assign m_1598_io_x1 = m_1183_io_cout; // @[MUL.scala 253:22]
  assign m_1598_io_x2 = m_1190_io_s; // @[MUL.scala 252:21]
  assign m_1598_io_x3 = m_1184_io_cout; // @[MUL.scala 253:22]
  assign m_1599_io_x1 = m_1191_io_s; // @[MUL.scala 252:21]
  assign m_1599_io_x2 = m_1185_io_cout; // @[MUL.scala 253:22]
  assign m_1599_io_x3 = m_1192_io_s; // @[MUL.scala 252:21]
  assign m_1600_io_x1 = m_1186_io_cout; // @[MUL.scala 253:22]
  assign m_1600_io_x2 = m_602_io_cout; // @[MUL.scala 253:22]
  assign m_1600_io_x3 = m_1187_io_out_1; // @[MUL.scala 105:13]
  assign m_1601_io_x1 = m_1193_io_s; // @[MUL.scala 252:21]
  assign m_1601_io_x2 = m_1188_io_cout; // @[MUL.scala 253:22]
  assign m_1601_io_x3 = m_1194_io_s; // @[MUL.scala 252:21]
  assign m_1602_io_x1 = m_1189_io_cout; // @[MUL.scala 253:22]
  assign m_1602_io_x2 = m_1195_io_s; // @[MUL.scala 252:21]
  assign m_1602_io_x3 = m_1190_io_cout; // @[MUL.scala 253:22]
  assign m_1603_io_x1 = m_1196_io_s; // @[MUL.scala 252:21]
  assign m_1603_io_x2 = m_1191_io_cout; // @[MUL.scala 253:22]
  assign m_1603_io_x3 = m_1197_io_s; // @[MUL.scala 252:21]
  assign m_1604_io_in_0 = m_1192_io_cout; // @[MUL.scala 253:22]
  assign m_1604_io_in_1 = m_610_io_cout; // @[MUL.scala 253:22]
  assign m_1605_io_x1 = m_1198_io_s; // @[MUL.scala 252:21]
  assign m_1605_io_x2 = m_1193_io_cout; // @[MUL.scala 253:22]
  assign m_1605_io_x3 = m_1199_io_s; // @[MUL.scala 252:21]
  assign m_1606_io_x1 = m_1194_io_cout; // @[MUL.scala 253:22]
  assign m_1606_io_x2 = m_1200_io_s; // @[MUL.scala 252:21]
  assign m_1606_io_x3 = m_1195_io_cout; // @[MUL.scala 253:22]
  assign m_1607_io_x1 = m_1201_io_s; // @[MUL.scala 252:21]
  assign m_1607_io_x2 = m_1196_io_cout; // @[MUL.scala 253:22]
  assign m_1607_io_x3 = m_1202_io_s; // @[MUL.scala 252:21]
  assign m_1608_io_in_0 = m_1197_io_cout; // @[MUL.scala 253:22]
  assign m_1608_io_in_1 = m_618_io_cout; // @[MUL.scala 253:22]
  assign m_1609_io_x1 = m_1203_io_s; // @[MUL.scala 252:21]
  assign m_1609_io_x2 = m_1198_io_cout; // @[MUL.scala 253:22]
  assign m_1609_io_x3 = m_1204_io_s; // @[MUL.scala 252:21]
  assign m_1610_io_x1 = m_1199_io_cout; // @[MUL.scala 253:22]
  assign m_1610_io_x2 = m_1205_io_s; // @[MUL.scala 252:21]
  assign m_1610_io_x3 = m_1200_io_cout; // @[MUL.scala 253:22]
  assign m_1611_io_x1 = m_1206_io_s; // @[MUL.scala 252:21]
  assign m_1611_io_x2 = m_1201_io_cout; // @[MUL.scala 253:22]
  assign m_1611_io_x3 = m_1207_io_s; // @[MUL.scala 252:21]
  assign m_1612_io_in_0 = m_1202_io_cout; // @[MUL.scala 253:22]
  assign m_1612_io_in_1 = m_626_io_out_1; // @[MUL.scala 126:16]
  assign m_1613_io_x1 = m_1208_io_s; // @[MUL.scala 252:21]
  assign m_1613_io_x2 = m_1203_io_cout; // @[MUL.scala 253:22]
  assign m_1613_io_x3 = m_1209_io_s; // @[MUL.scala 252:21]
  assign m_1614_io_x1 = m_1204_io_cout; // @[MUL.scala 253:22]
  assign m_1614_io_x2 = m_1210_io_s; // @[MUL.scala 252:21]
  assign m_1614_io_x3 = m_1205_io_cout; // @[MUL.scala 253:22]
  assign m_1615_io_x1 = m_1211_io_s; // @[MUL.scala 252:21]
  assign m_1615_io_x2 = m_1206_io_cout; // @[MUL.scala 253:22]
  assign m_1615_io_x3 = m_1212_io_s; // @[MUL.scala 252:21]
  assign m_1616_io_in_0 = m_1207_io_cout; // @[MUL.scala 253:22]
  assign m_1616_io_in_1 = m_634_io_out_1; // @[MUL.scala 126:16]
  assign m_1617_io_x1 = m_1213_io_s; // @[MUL.scala 252:21]
  assign m_1617_io_x2 = m_1208_io_cout; // @[MUL.scala 253:22]
  assign m_1617_io_x3 = m_1214_io_s; // @[MUL.scala 252:21]
  assign m_1618_io_x1 = m_1209_io_cout; // @[MUL.scala 253:22]
  assign m_1618_io_x2 = m_1215_io_s; // @[MUL.scala 252:21]
  assign m_1618_io_x3 = m_1210_io_cout; // @[MUL.scala 253:22]
  assign m_1619_io_x1 = m_1216_io_s; // @[MUL.scala 252:21]
  assign m_1619_io_x2 = m_1211_io_cout; // @[MUL.scala 253:22]
  assign m_1619_io_x3 = m_1217_io_s; // @[MUL.scala 252:21]
  assign m_1620_io_x1 = m_1218_io_s; // @[MUL.scala 252:21]
  assign m_1620_io_x2 = m_1213_io_cout; // @[MUL.scala 253:22]
  assign m_1620_io_x3 = m_1219_io_s; // @[MUL.scala 252:21]
  assign m_1621_io_x1 = m_1214_io_cout; // @[MUL.scala 253:22]
  assign m_1621_io_x2 = m_1220_io_s; // @[MUL.scala 252:21]
  assign m_1621_io_x3 = m_1215_io_cout; // @[MUL.scala 253:22]
  assign m_1622_io_x1 = m_1221_io_s; // @[MUL.scala 252:21]
  assign m_1622_io_x2 = m_1216_io_cout; // @[MUL.scala 253:22]
  assign m_1622_io_x3 = m_1222_io_out_0; // @[MUL.scala 105:13]
  assign m_1623_io_x1 = m_1223_io_s; // @[MUL.scala 252:21]
  assign m_1623_io_x2 = m_1218_io_cout; // @[MUL.scala 253:22]
  assign m_1623_io_x3 = m_1224_io_s; // @[MUL.scala 252:21]
  assign m_1624_io_x1 = m_1219_io_cout; // @[MUL.scala 253:22]
  assign m_1624_io_x2 = m_1225_io_s; // @[MUL.scala 252:21]
  assign m_1624_io_x3 = m_1220_io_cout; // @[MUL.scala 253:22]
  assign m_1625_io_x1 = m_1226_io_s; // @[MUL.scala 252:21]
  assign m_1625_io_x2 = m_1221_io_cout; // @[MUL.scala 253:22]
  assign m_1625_io_x3 = m_1227_io_out_0; // @[MUL.scala 105:13]
  assign m_1626_io_x1 = m_1228_io_s; // @[MUL.scala 252:21]
  assign m_1626_io_x2 = m_1223_io_cout; // @[MUL.scala 253:22]
  assign m_1626_io_x3 = m_1229_io_s; // @[MUL.scala 252:21]
  assign m_1627_io_x1 = m_1224_io_cout; // @[MUL.scala 253:22]
  assign m_1627_io_x2 = m_1230_io_s; // @[MUL.scala 252:21]
  assign m_1627_io_x3 = m_1225_io_cout; // @[MUL.scala 253:22]
  assign m_1628_io_x1 = m_1231_io_s; // @[MUL.scala 252:21]
  assign m_1628_io_x2 = m_1226_io_cout; // @[MUL.scala 253:22]
  assign m_1628_io_x3 = m_1232_io_out_0; // @[MUL.scala 105:13]
  assign m_1629_io_x1 = m_1233_io_s; // @[MUL.scala 252:21]
  assign m_1629_io_x2 = m_1228_io_cout; // @[MUL.scala 253:22]
  assign m_1629_io_x3 = m_1234_io_s; // @[MUL.scala 252:21]
  assign m_1630_io_x1 = m_1229_io_cout; // @[MUL.scala 253:22]
  assign m_1630_io_x2 = m_1235_io_s; // @[MUL.scala 252:21]
  assign m_1630_io_x3 = m_1230_io_cout; // @[MUL.scala 253:22]
  assign m_1631_io_x1 = m_1236_io_s; // @[MUL.scala 252:21]
  assign m_1631_io_x2 = m_1231_io_cout; // @[MUL.scala 253:22]
  assign m_1631_io_x3 = m_1237_io_out_0; // @[MUL.scala 105:13]
  assign m_1632_io_x1 = m_1238_io_s; // @[MUL.scala 252:21]
  assign m_1632_io_x2 = m_1233_io_cout; // @[MUL.scala 253:22]
  assign m_1632_io_x3 = m_1239_io_s; // @[MUL.scala 252:21]
  assign m_1633_io_x1 = m_1234_io_cout; // @[MUL.scala 253:22]
  assign m_1633_io_x2 = m_1240_io_s; // @[MUL.scala 252:21]
  assign m_1633_io_x3 = m_1235_io_cout; // @[MUL.scala 253:22]
  assign m_1634_io_x1 = m_1241_io_s; // @[MUL.scala 252:21]
  assign m_1634_io_x2 = m_1236_io_cout; // @[MUL.scala 253:22]
  assign m_1634_io_x3 = m_1242_io_out_0; // @[MUL.scala 105:13]
  assign m_1635_io_x1 = m_1243_io_s; // @[MUL.scala 252:21]
  assign m_1635_io_x2 = m_1238_io_cout; // @[MUL.scala 253:22]
  assign m_1635_io_x3 = m_1244_io_s; // @[MUL.scala 252:21]
  assign m_1636_io_x1 = m_1239_io_cout; // @[MUL.scala 253:22]
  assign m_1636_io_x2 = m_1245_io_s; // @[MUL.scala 252:21]
  assign m_1636_io_x3 = m_1240_io_cout; // @[MUL.scala 253:22]
  assign m_1637_io_x1 = m_1246_io_s; // @[MUL.scala 252:21]
  assign m_1637_io_x2 = m_1241_io_cout; // @[MUL.scala 253:22]
  assign m_1637_io_x3 = r_1966; // @[MUL.scala 105:13]
  assign m_1638_io_x1 = m_1247_io_s; // @[MUL.scala 252:21]
  assign m_1638_io_x2 = m_1243_io_cout; // @[MUL.scala 253:22]
  assign m_1638_io_x3 = m_1248_io_s; // @[MUL.scala 252:21]
  assign m_1639_io_x1 = m_1244_io_cout; // @[MUL.scala 253:22]
  assign m_1639_io_x2 = m_1249_io_s; // @[MUL.scala 252:21]
  assign m_1639_io_x3 = m_1245_io_cout; // @[MUL.scala 253:22]
  assign m_1640_io_in_0 = m_1250_io_s; // @[MUL.scala 252:21]
  assign m_1640_io_in_1 = m_1246_io_cout; // @[MUL.scala 253:22]
  assign m_1641_io_x1 = m_1251_io_s; // @[MUL.scala 252:21]
  assign m_1641_io_x2 = m_1247_io_cout; // @[MUL.scala 253:22]
  assign m_1641_io_x3 = m_1252_io_s; // @[MUL.scala 252:21]
  assign m_1642_io_x1 = m_1248_io_cout; // @[MUL.scala 253:22]
  assign m_1642_io_x2 = m_1253_io_s; // @[MUL.scala 252:21]
  assign m_1642_io_x3 = m_1249_io_cout; // @[MUL.scala 253:22]
  assign m_1643_io_in_0 = m_1254_io_s; // @[MUL.scala 252:21]
  assign m_1643_io_in_1 = m_1250_io_cout; // @[MUL.scala 253:22]
  assign m_1644_io_x1 = m_1255_io_s; // @[MUL.scala 252:21]
  assign m_1644_io_x2 = m_1251_io_cout; // @[MUL.scala 253:22]
  assign m_1644_io_x3 = m_1256_io_s; // @[MUL.scala 252:21]
  assign m_1645_io_x1 = m_1252_io_cout; // @[MUL.scala 253:22]
  assign m_1645_io_x2 = m_1257_io_s; // @[MUL.scala 252:21]
  assign m_1645_io_x3 = m_1253_io_cout; // @[MUL.scala 253:22]
  assign m_1646_io_in_0 = m_1258_io_s; // @[MUL.scala 252:21]
  assign m_1646_io_in_1 = m_1254_io_cout; // @[MUL.scala 253:22]
  assign m_1647_io_x1 = m_1259_io_s; // @[MUL.scala 252:21]
  assign m_1647_io_x2 = m_1255_io_cout; // @[MUL.scala 253:22]
  assign m_1647_io_x3 = m_1260_io_s; // @[MUL.scala 252:21]
  assign m_1648_io_x1 = m_1256_io_cout; // @[MUL.scala 253:22]
  assign m_1648_io_x2 = m_1261_io_s; // @[MUL.scala 252:21]
  assign m_1648_io_x3 = m_1257_io_cout; // @[MUL.scala 253:22]
  assign m_1649_io_in_0 = m_1262_io_s; // @[MUL.scala 252:21]
  assign m_1649_io_in_1 = m_1258_io_cout; // @[MUL.scala 253:22]
  assign m_1650_io_x1 = m_1263_io_s; // @[MUL.scala 252:21]
  assign m_1650_io_x2 = m_1259_io_cout; // @[MUL.scala 253:22]
  assign m_1650_io_x3 = m_1264_io_s; // @[MUL.scala 252:21]
  assign m_1651_io_x1 = m_1260_io_cout; // @[MUL.scala 253:22]
  assign m_1651_io_x2 = m_1265_io_s; // @[MUL.scala 252:21]
  assign m_1651_io_x3 = m_1261_io_cout; // @[MUL.scala 253:22]
  assign m_1652_io_in_0 = m_1266_io_s; // @[MUL.scala 252:21]
  assign m_1652_io_in_1 = m_1262_io_cout; // @[MUL.scala 253:22]
  assign m_1653_io_x1 = m_1267_io_s; // @[MUL.scala 252:21]
  assign m_1653_io_x2 = m_1263_io_cout; // @[MUL.scala 253:22]
  assign m_1653_io_x3 = m_1268_io_s; // @[MUL.scala 252:21]
  assign m_1654_io_x1 = m_1264_io_cout; // @[MUL.scala 253:22]
  assign m_1654_io_x2 = m_1269_io_s; // @[MUL.scala 252:21]
  assign m_1654_io_x3 = m_1265_io_cout; // @[MUL.scala 253:22]
  assign m_1655_io_in_0 = m_1270_io_out_0; // @[MUL.scala 125:16]
  assign m_1655_io_in_1 = m_1266_io_cout; // @[MUL.scala 253:22]
  assign m_1656_io_x1 = m_1271_io_s; // @[MUL.scala 252:21]
  assign m_1656_io_x2 = m_1267_io_cout; // @[MUL.scala 253:22]
  assign m_1656_io_x3 = m_1272_io_s; // @[MUL.scala 252:21]
  assign m_1657_io_x1 = m_1268_io_cout; // @[MUL.scala 253:22]
  assign m_1657_io_x2 = m_1273_io_s; // @[MUL.scala 252:21]
  assign m_1657_io_x3 = m_1269_io_cout; // @[MUL.scala 253:22]
  assign m_1658_io_in_0 = m_722_io_cout; // @[MUL.scala 253:22]
  assign m_1658_io_in_1 = m_1270_io_out_1; // @[MUL.scala 126:16]
  assign m_1659_io_x1 = m_1274_io_s; // @[MUL.scala 252:21]
  assign m_1659_io_x2 = m_1271_io_cout; // @[MUL.scala 253:22]
  assign m_1659_io_x3 = m_1275_io_s; // @[MUL.scala 252:21]
  assign m_1660_io_x1 = m_1272_io_cout; // @[MUL.scala 253:22]
  assign m_1660_io_x2 = m_1276_io_s; // @[MUL.scala 252:21]
  assign m_1660_io_x3 = m_1273_io_cout; // @[MUL.scala 253:22]
  assign m_1661_io_x1 = m_1277_io_s; // @[MUL.scala 252:21]
  assign m_1661_io_x2 = m_1274_io_cout; // @[MUL.scala 253:22]
  assign m_1661_io_x3 = m_1278_io_s; // @[MUL.scala 252:21]
  assign m_1662_io_x1 = m_1275_io_cout; // @[MUL.scala 253:22]
  assign m_1662_io_x2 = m_1279_io_s; // @[MUL.scala 252:21]
  assign m_1662_io_x3 = m_1276_io_cout; // @[MUL.scala 253:22]
  assign m_1663_io_x1 = m_1280_io_s; // @[MUL.scala 252:21]
  assign m_1663_io_x2 = m_1277_io_cout; // @[MUL.scala 253:22]
  assign m_1663_io_x3 = m_1281_io_s; // @[MUL.scala 252:21]
  assign m_1664_io_x1 = m_1278_io_cout; // @[MUL.scala 253:22]
  assign m_1664_io_x2 = m_1282_io_s; // @[MUL.scala 252:21]
  assign m_1664_io_x3 = m_1279_io_cout; // @[MUL.scala 253:22]
  assign m_1665_io_x1 = m_1283_io_s; // @[MUL.scala 252:21]
  assign m_1665_io_x2 = m_1280_io_cout; // @[MUL.scala 253:22]
  assign m_1665_io_x3 = m_1284_io_s; // @[MUL.scala 252:21]
  assign m_1666_io_x1 = m_1281_io_cout; // @[MUL.scala 253:22]
  assign m_1666_io_x2 = m_1285_io_s; // @[MUL.scala 252:21]
  assign m_1666_io_x3 = m_1282_io_cout; // @[MUL.scala 253:22]
  assign m_1667_io_x1 = m_1286_io_s; // @[MUL.scala 252:21]
  assign m_1667_io_x2 = m_1283_io_cout; // @[MUL.scala 253:22]
  assign m_1667_io_x3 = m_1287_io_s; // @[MUL.scala 252:21]
  assign m_1668_io_x1 = m_1284_io_cout; // @[MUL.scala 253:22]
  assign m_1668_io_x2 = m_1288_io_s; // @[MUL.scala 252:21]
  assign m_1668_io_x3 = m_1285_io_cout; // @[MUL.scala 253:22]
  assign m_1669_io_x1 = m_1289_io_s; // @[MUL.scala 252:21]
  assign m_1669_io_x2 = m_1286_io_cout; // @[MUL.scala 253:22]
  assign m_1669_io_x3 = m_1290_io_s; // @[MUL.scala 252:21]
  assign m_1670_io_x1 = m_1287_io_cout; // @[MUL.scala 253:22]
  assign m_1670_io_x2 = m_1291_io_out_0; // @[MUL.scala 104:13]
  assign m_1670_io_x3 = m_1288_io_cout; // @[MUL.scala 253:22]
  assign m_1671_io_x1 = m_1292_io_s; // @[MUL.scala 252:21]
  assign m_1671_io_x2 = m_1289_io_cout; // @[MUL.scala 253:22]
  assign m_1671_io_x3 = m_1293_io_s; // @[MUL.scala 252:21]
  assign m_1672_io_x1 = m_1290_io_cout; // @[MUL.scala 253:22]
  assign m_1672_io_x2 = m_1294_io_out_0; // @[MUL.scala 104:13]
  assign m_1672_io_x3 = m_1291_io_out_1; // @[MUL.scala 105:13]
  assign m_1673_io_x1 = m_1295_io_s; // @[MUL.scala 252:21]
  assign m_1673_io_x2 = m_1292_io_cout; // @[MUL.scala 253:22]
  assign m_1673_io_x3 = m_1296_io_s; // @[MUL.scala 252:21]
  assign m_1674_io_x1 = m_1293_io_cout; // @[MUL.scala 253:22]
  assign m_1674_io_x2 = m_1297_io_out_0; // @[MUL.scala 104:13]
  assign m_1674_io_x3 = m_1294_io_out_1; // @[MUL.scala 105:13]
  assign m_1675_io_x1 = m_1298_io_s; // @[MUL.scala 252:21]
  assign m_1675_io_x2 = m_1295_io_cout; // @[MUL.scala 253:22]
  assign m_1675_io_x3 = m_1299_io_s; // @[MUL.scala 252:21]
  assign m_1676_io_x1 = m_1296_io_cout; // @[MUL.scala 253:22]
  assign m_1676_io_x2 = m_1300_io_out_0; // @[MUL.scala 104:13]
  assign m_1676_io_x3 = m_1297_io_out_1; // @[MUL.scala 105:13]
  assign m_1677_io_x1 = m_1301_io_s; // @[MUL.scala 252:21]
  assign m_1677_io_x2 = m_1298_io_cout; // @[MUL.scala 253:22]
  assign m_1677_io_x3 = m_1302_io_s; // @[MUL.scala 252:21]
  assign m_1678_io_x1 = m_1299_io_cout; // @[MUL.scala 253:22]
  assign m_1678_io_x2 = m_1303_io_out_0; // @[MUL.scala 104:13]
  assign m_1678_io_x3 = m_1300_io_out_1; // @[MUL.scala 105:13]
  assign m_1679_io_x1 = m_1304_io_s; // @[MUL.scala 252:21]
  assign m_1679_io_x2 = m_1301_io_cout; // @[MUL.scala 253:22]
  assign m_1679_io_x3 = m_1305_io_s; // @[MUL.scala 252:21]
  assign m_1680_io_x1 = m_1302_io_cout; // @[MUL.scala 253:22]
  assign m_1680_io_x2 = r_2218; // @[MUL.scala 104:13]
  assign m_1680_io_x3 = m_1303_io_out_1; // @[MUL.scala 105:13]
  assign m_1681_io_x1 = m_1306_io_s; // @[MUL.scala 252:21]
  assign m_1681_io_x2 = m_1304_io_cout; // @[MUL.scala 253:22]
  assign m_1681_io_x3 = m_1307_io_s; // @[MUL.scala 252:21]
  assign m_1682_io_x1 = m_1308_io_s; // @[MUL.scala 252:21]
  assign m_1682_io_x2 = m_1306_io_cout; // @[MUL.scala 253:22]
  assign m_1682_io_x3 = m_1309_io_s; // @[MUL.scala 252:21]
  assign m_1683_io_x1 = m_1310_io_s; // @[MUL.scala 252:21]
  assign m_1683_io_x2 = m_1308_io_cout; // @[MUL.scala 253:22]
  assign m_1683_io_x3 = m_1311_io_s; // @[MUL.scala 252:21]
  assign m_1684_io_x1 = m_1312_io_s; // @[MUL.scala 252:21]
  assign m_1684_io_x2 = m_1310_io_cout; // @[MUL.scala 253:22]
  assign m_1684_io_x3 = m_1313_io_s; // @[MUL.scala 252:21]
  assign m_1685_io_x1 = m_1314_io_s; // @[MUL.scala 252:21]
  assign m_1685_io_x2 = m_1312_io_cout; // @[MUL.scala 253:22]
  assign m_1685_io_x3 = m_1315_io_s; // @[MUL.scala 252:21]
  assign m_1686_io_x1 = m_1316_io_s; // @[MUL.scala 252:21]
  assign m_1686_io_x2 = m_1314_io_cout; // @[MUL.scala 253:22]
  assign m_1686_io_x3 = m_1317_io_out_0; // @[MUL.scala 105:13]
  assign m_1687_io_x1 = m_1318_io_s; // @[MUL.scala 252:21]
  assign m_1687_io_x2 = m_1316_io_cout; // @[MUL.scala 253:22]
  assign m_1687_io_x3 = m_788_io_cout; // @[MUL.scala 253:22]
  assign m_1688_io_x1 = m_1319_io_s; // @[MUL.scala 252:21]
  assign m_1688_io_x2 = m_1318_io_cout; // @[MUL.scala 253:22]
  assign m_1688_io_x3 = m_790_io_cout; // @[MUL.scala 253:22]
  assign m_1689_io_x1 = m_1320_io_s; // @[MUL.scala 252:21]
  assign m_1689_io_x2 = m_1319_io_cout; // @[MUL.scala 253:22]
  assign m_1689_io_x3 = m_792_io_cout; // @[MUL.scala 253:22]
  assign m_1690_io_x1 = m_1321_io_s; // @[MUL.scala 252:21]
  assign m_1690_io_x2 = m_1320_io_cout; // @[MUL.scala 253:22]
  assign m_1690_io_x3 = m_794_io_out_1; // @[MUL.scala 105:13]
  assign m_1691_io_x1 = m_1322_io_s; // @[MUL.scala 252:21]
  assign m_1691_io_x2 = m_1321_io_cout; // @[MUL.scala 253:22]
  assign m_1691_io_x3 = m_796_io_out_1; // @[MUL.scala 105:13]
  assign m_1692_io_in_0 = m_1323_io_s; // @[MUL.scala 252:21]
  assign m_1692_io_in_1 = m_1322_io_cout; // @[MUL.scala 253:22]
  assign m_1693_io_in_0 = m_1324_io_out_0; // @[MUL.scala 125:16]
  assign m_1693_io_in_1 = m_1323_io_cout; // @[MUL.scala 253:22]
  assign m_1694_io_in_0 = m_1325_io_out_0; // @[MUL.scala 125:16]
  assign m_1694_io_in_1 = m_1324_io_out_1; // @[MUL.scala 126:16]
  assign m_1695_io_in_0 = m_1326_io_out_0; // @[MUL.scala 125:16]
  assign m_1695_io_in_1 = m_1325_io_out_1; // @[MUL.scala 126:16]
  assign m_1696_io_in_0 = m_1327_io_out_0; // @[MUL.scala 125:16]
  assign m_1696_io_in_1 = m_1326_io_out_1; // @[MUL.scala 126:16]
  assign m_1697_io_in_0 = m_1328_io_out_0; // @[MUL.scala 125:16]
  assign m_1697_io_in_1 = m_1327_io_out_1; // @[MUL.scala 126:16]
  assign m_1698_io_in_0 = m_1330_io_out_0; // @[MUL.scala 125:16]
  assign m_1698_io_in_1 = m_1329_io_out_1; // @[MUL.scala 126:16]
  assign m_1699_io_in_0 = m_1331_io_out_0; // @[MUL.scala 125:16]
  assign m_1699_io_in_1 = m_1330_io_out_1; // @[MUL.scala 126:16]
  assign m_1700_io_in_0 = m_1332_io_out_0; // @[MUL.scala 125:16]
  assign m_1700_io_in_1 = m_1331_io_out_1; // @[MUL.scala 126:16]
  assign m_1701_io_in_0 = m_1333_io_out_0; // @[MUL.scala 125:16]
  assign m_1701_io_in_1 = m_1332_io_out_1; // @[MUL.scala 126:16]
  assign m_1702_io_in_0 = m_1334_io_s; // @[MUL.scala 252:21]
  assign m_1702_io_in_1 = m_1333_io_out_1; // @[MUL.scala 126:16]
  assign m_1703_io_in_0 = m_1335_io_s; // @[MUL.scala 252:21]
  assign m_1703_io_in_1 = m_1334_io_cout; // @[MUL.scala 253:22]
  assign m_1704_io_in_0 = m_1336_io_s; // @[MUL.scala 252:21]
  assign m_1704_io_in_1 = m_1335_io_cout; // @[MUL.scala 253:22]
  assign m_1705_io_in_0 = m_1337_io_s; // @[MUL.scala 252:21]
  assign m_1705_io_in_1 = m_1336_io_cout; // @[MUL.scala 253:22]
  assign m_1706_io_x1 = m_1338_io_s; // @[MUL.scala 252:21]
  assign m_1706_io_x2 = m_1337_io_cout; // @[MUL.scala 253:22]
  assign m_1706_io_x3 = m_813_io_out_1; // @[MUL.scala 105:13]
  assign m_1707_io_x1 = m_1339_io_s; // @[MUL.scala 252:21]
  assign m_1707_io_x2 = m_1338_io_cout; // @[MUL.scala 253:22]
  assign m_1707_io_x3 = m_815_io_out_1; // @[MUL.scala 105:13]
  assign m_1708_io_x1 = m_1340_io_s; // @[MUL.scala 252:21]
  assign m_1708_io_x2 = m_1339_io_cout; // @[MUL.scala 253:22]
  assign m_1708_io_x3 = m_817_io_out_1; // @[MUL.scala 105:13]
  assign m_1709_io_x1 = m_1341_io_s; // @[MUL.scala 252:21]
  assign m_1709_io_x2 = m_1340_io_cout; // @[MUL.scala 253:22]
  assign m_1709_io_x3 = m_819_io_cout; // @[MUL.scala 253:22]
  assign m_1710_io_x1 = m_1342_io_s; // @[MUL.scala 252:21]
  assign m_1710_io_x2 = m_1341_io_cout; // @[MUL.scala 253:22]
  assign m_1710_io_x3 = m_821_io_cout; // @[MUL.scala 253:22]
  assign m_1711_io_x1 = m_1343_io_s; // @[MUL.scala 252:21]
  assign m_1711_io_x2 = m_1342_io_cout; // @[MUL.scala 253:22]
  assign m_1711_io_x3 = m_1344_io_out_0; // @[MUL.scala 105:13]
  assign m_1712_io_x1 = m_1345_io_s; // @[MUL.scala 252:21]
  assign m_1712_io_x2 = m_1343_io_cout; // @[MUL.scala 253:22]
  assign m_1712_io_x3 = m_1346_io_out_0; // @[MUL.scala 105:13]
  assign m_1713_io_x1 = m_1347_io_s; // @[MUL.scala 252:21]
  assign m_1713_io_x2 = m_1345_io_cout; // @[MUL.scala 253:22]
  assign m_1713_io_x3 = m_1348_io_out_0; // @[MUL.scala 105:13]
  assign m_1714_io_x1 = m_1349_io_s; // @[MUL.scala 252:21]
  assign m_1714_io_x2 = m_1347_io_cout; // @[MUL.scala 253:22]
  assign m_1714_io_x3 = m_1350_io_out_0; // @[MUL.scala 105:13]
  assign m_1715_io_x1 = m_1351_io_s; // @[MUL.scala 252:21]
  assign m_1715_io_x2 = m_1349_io_cout; // @[MUL.scala 253:22]
  assign m_1715_io_x3 = m_1352_io_s; // @[MUL.scala 252:21]
  assign m_1716_io_x1 = m_1353_io_s; // @[MUL.scala 252:21]
  assign m_1716_io_x2 = m_1351_io_cout; // @[MUL.scala 253:22]
  assign m_1716_io_x3 = m_1354_io_s; // @[MUL.scala 252:21]
  assign m_1717_io_x1 = m_1355_io_s; // @[MUL.scala 252:21]
  assign m_1717_io_x2 = m_1353_io_cout; // @[MUL.scala 253:22]
  assign m_1717_io_x3 = m_1356_io_s; // @[MUL.scala 252:21]
  assign m_1718_io_x1 = m_1357_io_s; // @[MUL.scala 252:21]
  assign m_1718_io_x2 = m_1355_io_cout; // @[MUL.scala 253:22]
  assign m_1718_io_x3 = m_1358_io_s; // @[MUL.scala 252:21]
  assign m_1719_io_x1 = m_1359_io_s; // @[MUL.scala 252:21]
  assign m_1719_io_x2 = m_1357_io_cout; // @[MUL.scala 253:22]
  assign m_1719_io_x3 = m_1360_io_s; // @[MUL.scala 252:21]
  assign m_1720_io_x1 = m_1361_io_s; // @[MUL.scala 252:21]
  assign m_1720_io_x2 = m_1359_io_cout; // @[MUL.scala 253:22]
  assign m_1720_io_x3 = m_1362_io_s; // @[MUL.scala 252:21]
  assign m_1721_io_in_0 = m_1360_io_cout; // @[MUL.scala 253:22]
  assign m_1721_io_in_1 = m_97_io_out_1; // @[MUL.scala 126:16]
  assign m_1722_io_x1 = m_1363_io_s; // @[MUL.scala 252:21]
  assign m_1722_io_x2 = m_1361_io_cout; // @[MUL.scala 253:22]
  assign m_1722_io_x3 = m_1364_io_s; // @[MUL.scala 252:21]
  assign m_1723_io_in_0 = m_1362_io_cout; // @[MUL.scala 253:22]
  assign m_1723_io_in_1 = m_102_io_out_1; // @[MUL.scala 126:16]
  assign m_1724_io_x1 = m_1365_io_s; // @[MUL.scala 252:21]
  assign m_1724_io_x2 = m_1363_io_cout; // @[MUL.scala 253:22]
  assign m_1724_io_x3 = m_1366_io_s; // @[MUL.scala 252:21]
  assign m_1725_io_in_0 = m_1364_io_cout; // @[MUL.scala 253:22]
  assign m_1725_io_in_1 = m_107_io_cout; // @[MUL.scala 253:22]
  assign m_1726_io_x1 = m_1367_io_s; // @[MUL.scala 252:21]
  assign m_1726_io_x2 = m_1365_io_cout; // @[MUL.scala 253:22]
  assign m_1726_io_x3 = m_1368_io_s; // @[MUL.scala 252:21]
  assign m_1727_io_in_0 = m_1366_io_cout; // @[MUL.scala 253:22]
  assign m_1727_io_in_1 = m_860_io_out_0; // @[MUL.scala 126:16]
  assign m_1728_io_x1 = m_1369_io_s; // @[MUL.scala 252:21]
  assign m_1728_io_x2 = m_1367_io_cout; // @[MUL.scala 253:22]
  assign m_1728_io_x3 = m_1370_io_s; // @[MUL.scala 252:21]
  assign m_1729_io_in_0 = m_1368_io_cout; // @[MUL.scala 253:22]
  assign m_1729_io_in_1 = m_1371_io_out_0; // @[MUL.scala 126:16]
  assign m_1730_io_x1 = m_1372_io_s; // @[MUL.scala 252:21]
  assign m_1730_io_x2 = m_1369_io_cout; // @[MUL.scala 253:22]
  assign m_1730_io_x3 = m_1373_io_s; // @[MUL.scala 252:21]
  assign m_1731_io_x1 = m_1370_io_cout; // @[MUL.scala 253:22]
  assign m_1731_io_x2 = m_1374_io_out_0; // @[MUL.scala 104:13]
  assign m_1731_io_x3 = m_1371_io_out_1; // @[MUL.scala 105:13]
  assign m_1732_io_x1 = m_1375_io_s; // @[MUL.scala 252:21]
  assign m_1732_io_x2 = m_1372_io_cout; // @[MUL.scala 253:22]
  assign m_1732_io_x3 = m_1376_io_s; // @[MUL.scala 252:21]
  assign m_1733_io_x1 = m_1373_io_cout; // @[MUL.scala 253:22]
  assign m_1733_io_x2 = m_1377_io_out_0; // @[MUL.scala 104:13]
  assign m_1733_io_x3 = m_1374_io_out_1; // @[MUL.scala 105:13]
  assign m_1734_io_x1 = m_1378_io_s; // @[MUL.scala 252:21]
  assign m_1734_io_x2 = m_1375_io_cout; // @[MUL.scala 253:22]
  assign m_1734_io_x3 = m_1379_io_s; // @[MUL.scala 252:21]
  assign m_1735_io_x1 = m_1376_io_cout; // @[MUL.scala 253:22]
  assign m_1735_io_x2 = m_1380_io_out_0; // @[MUL.scala 104:13]
  assign m_1735_io_x3 = m_1377_io_out_1; // @[MUL.scala 105:13]
  assign m_1736_io_x1 = m_1381_io_s; // @[MUL.scala 252:21]
  assign m_1736_io_x2 = m_1378_io_cout; // @[MUL.scala 253:22]
  assign m_1736_io_x3 = m_1382_io_s; // @[MUL.scala 252:21]
  assign m_1737_io_x1 = m_1379_io_cout; // @[MUL.scala 253:22]
  assign m_1737_io_x2 = m_1383_io_out_0; // @[MUL.scala 104:13]
  assign m_1737_io_x3 = m_1380_io_out_1; // @[MUL.scala 105:13]
  assign m_1738_io_x1 = m_1384_io_s; // @[MUL.scala 252:21]
  assign m_1738_io_x2 = m_1381_io_cout; // @[MUL.scala 253:22]
  assign m_1738_io_x3 = m_1385_io_s; // @[MUL.scala 252:21]
  assign m_1739_io_x1 = m_1382_io_cout; // @[MUL.scala 253:22]
  assign m_1739_io_x2 = m_1386_io_s; // @[MUL.scala 252:21]
  assign m_1739_io_x3 = m_1383_io_out_1; // @[MUL.scala 105:13]
  assign m_1740_io_x1 = m_1387_io_s; // @[MUL.scala 252:21]
  assign m_1740_io_x2 = m_1384_io_cout; // @[MUL.scala 253:22]
  assign m_1740_io_x3 = m_1388_io_s; // @[MUL.scala 252:21]
  assign m_1741_io_x1 = m_1385_io_cout; // @[MUL.scala 253:22]
  assign m_1741_io_x2 = m_1389_io_s; // @[MUL.scala 252:21]
  assign m_1741_io_x3 = m_1386_io_cout; // @[MUL.scala 253:22]
  assign m_1742_io_x1 = m_1390_io_s; // @[MUL.scala 252:21]
  assign m_1742_io_x2 = m_1387_io_cout; // @[MUL.scala 253:22]
  assign m_1742_io_x3 = m_1391_io_s; // @[MUL.scala 252:21]
  assign m_1743_io_x1 = m_1388_io_cout; // @[MUL.scala 253:22]
  assign m_1743_io_x2 = m_1392_io_s; // @[MUL.scala 252:21]
  assign m_1743_io_x3 = m_1389_io_cout; // @[MUL.scala 253:22]
  assign m_1744_io_x1 = m_1393_io_s; // @[MUL.scala 252:21]
  assign m_1744_io_x2 = m_1390_io_cout; // @[MUL.scala 253:22]
  assign m_1744_io_x3 = m_1394_io_s; // @[MUL.scala 252:21]
  assign m_1745_io_x1 = m_1391_io_cout; // @[MUL.scala 253:22]
  assign m_1745_io_x2 = m_1395_io_s; // @[MUL.scala 252:21]
  assign m_1745_io_x3 = m_1392_io_cout; // @[MUL.scala 253:22]
  assign m_1746_io_x1 = m_1396_io_s; // @[MUL.scala 252:21]
  assign m_1746_io_x2 = m_1393_io_cout; // @[MUL.scala 253:22]
  assign m_1746_io_x3 = m_1397_io_s; // @[MUL.scala 252:21]
  assign m_1747_io_x1 = m_1394_io_cout; // @[MUL.scala 253:22]
  assign m_1747_io_x2 = m_1398_io_s; // @[MUL.scala 252:21]
  assign m_1747_io_x3 = m_1395_io_cout; // @[MUL.scala 253:22]
  assign m_1748_io_x1 = m_1399_io_s; // @[MUL.scala 252:21]
  assign m_1748_io_x2 = m_1396_io_cout; // @[MUL.scala 253:22]
  assign m_1748_io_x3 = m_1400_io_s; // @[MUL.scala 252:21]
  assign m_1749_io_x1 = m_1397_io_cout; // @[MUL.scala 253:22]
  assign m_1749_io_x2 = m_1401_io_s; // @[MUL.scala 252:21]
  assign m_1749_io_x3 = m_1398_io_cout; // @[MUL.scala 253:22]
  assign m_1750_io_x1 = m_1402_io_s; // @[MUL.scala 252:21]
  assign m_1750_io_x2 = m_1399_io_cout; // @[MUL.scala 253:22]
  assign m_1750_io_x3 = m_1403_io_s; // @[MUL.scala 252:21]
  assign m_1751_io_x1 = m_1400_io_cout; // @[MUL.scala 253:22]
  assign m_1751_io_x2 = m_1404_io_s; // @[MUL.scala 252:21]
  assign m_1751_io_x3 = m_1401_io_cout; // @[MUL.scala 253:22]
  assign m_1752_io_x1 = m_1405_io_s; // @[MUL.scala 252:21]
  assign m_1752_io_x2 = m_1402_io_cout; // @[MUL.scala 253:22]
  assign m_1752_io_x3 = m_1406_io_s; // @[MUL.scala 252:21]
  assign m_1753_io_x1 = m_1403_io_cout; // @[MUL.scala 253:22]
  assign m_1753_io_x2 = m_1407_io_s; // @[MUL.scala 252:21]
  assign m_1753_io_x3 = m_1404_io_cout; // @[MUL.scala 253:22]
  assign m_1754_io_x1 = m_1408_io_s; // @[MUL.scala 252:21]
  assign m_1754_io_x2 = m_1405_io_cout; // @[MUL.scala 253:22]
  assign m_1754_io_x3 = m_1409_io_s; // @[MUL.scala 252:21]
  assign m_1755_io_x1 = m_1406_io_cout; // @[MUL.scala 253:22]
  assign m_1755_io_x2 = m_1410_io_s; // @[MUL.scala 252:21]
  assign m_1755_io_x3 = m_1407_io_cout; // @[MUL.scala 253:22]
  assign m_1756_io_x1 = m_1411_io_s; // @[MUL.scala 252:21]
  assign m_1756_io_x2 = m_1408_io_cout; // @[MUL.scala 253:22]
  assign m_1756_io_x3 = m_1412_io_s; // @[MUL.scala 252:21]
  assign m_1757_io_x1 = m_1409_io_cout; // @[MUL.scala 253:22]
  assign m_1757_io_x2 = m_1413_io_s; // @[MUL.scala 252:21]
  assign m_1757_io_x3 = m_1410_io_cout; // @[MUL.scala 253:22]
  assign m_1758_io_x1 = m_1415_io_s; // @[MUL.scala 252:21]
  assign m_1758_io_x2 = m_1411_io_cout; // @[MUL.scala 253:22]
  assign m_1758_io_x3 = m_1416_io_s; // @[MUL.scala 252:21]
  assign m_1759_io_x1 = m_1412_io_cout; // @[MUL.scala 253:22]
  assign m_1759_io_x2 = m_1417_io_s; // @[MUL.scala 252:21]
  assign m_1759_io_x3 = m_1413_io_cout; // @[MUL.scala 253:22]
  assign m_1760_io_in_0 = m_1418_io_out_0; // @[MUL.scala 125:16]
  assign m_1760_io_in_1 = m_1414_io_out_1; // @[MUL.scala 126:16]
  assign m_1761_io_x1 = m_1419_io_s; // @[MUL.scala 252:21]
  assign m_1761_io_x2 = m_1415_io_cout; // @[MUL.scala 253:22]
  assign m_1761_io_x3 = m_1420_io_s; // @[MUL.scala 252:21]
  assign m_1762_io_x1 = m_1416_io_cout; // @[MUL.scala 253:22]
  assign m_1762_io_x2 = m_1421_io_s; // @[MUL.scala 252:21]
  assign m_1762_io_x3 = m_1417_io_cout; // @[MUL.scala 253:22]
  assign m_1763_io_in_0 = m_1422_io_out_0; // @[MUL.scala 125:16]
  assign m_1763_io_in_1 = m_1418_io_out_1; // @[MUL.scala 126:16]
  assign m_1764_io_x1 = m_1423_io_s; // @[MUL.scala 252:21]
  assign m_1764_io_x2 = m_1419_io_cout; // @[MUL.scala 253:22]
  assign m_1764_io_x3 = m_1424_io_s; // @[MUL.scala 252:21]
  assign m_1765_io_x1 = m_1420_io_cout; // @[MUL.scala 253:22]
  assign m_1765_io_x2 = m_1425_io_s; // @[MUL.scala 252:21]
  assign m_1765_io_x3 = m_1421_io_cout; // @[MUL.scala 253:22]
  assign m_1766_io_in_0 = m_1426_io_out_0; // @[MUL.scala 125:16]
  assign m_1766_io_in_1 = m_1422_io_out_1; // @[MUL.scala 126:16]
  assign m_1767_io_x1 = m_1427_io_s; // @[MUL.scala 252:21]
  assign m_1767_io_x2 = m_1423_io_cout; // @[MUL.scala 253:22]
  assign m_1767_io_x3 = m_1428_io_s; // @[MUL.scala 252:21]
  assign m_1768_io_x1 = m_1424_io_cout; // @[MUL.scala 253:22]
  assign m_1768_io_x2 = m_1429_io_s; // @[MUL.scala 252:21]
  assign m_1768_io_x3 = m_1425_io_cout; // @[MUL.scala 253:22]
  assign m_1769_io_in_0 = m_1430_io_s; // @[MUL.scala 252:21]
  assign m_1769_io_in_1 = m_1426_io_out_1; // @[MUL.scala 126:16]
  assign m_1770_io_x1 = m_1431_io_s; // @[MUL.scala 252:21]
  assign m_1770_io_x2 = m_1427_io_cout; // @[MUL.scala 253:22]
  assign m_1770_io_x3 = m_1432_io_s; // @[MUL.scala 252:21]
  assign m_1771_io_x1 = m_1428_io_cout; // @[MUL.scala 253:22]
  assign m_1771_io_x2 = m_1433_io_s; // @[MUL.scala 252:21]
  assign m_1771_io_x3 = m_1429_io_cout; // @[MUL.scala 253:22]
  assign m_1772_io_in_0 = m_1434_io_s; // @[MUL.scala 252:21]
  assign m_1772_io_in_1 = m_1430_io_cout; // @[MUL.scala 253:22]
  assign m_1773_io_x1 = m_1435_io_s; // @[MUL.scala 252:21]
  assign m_1773_io_x2 = m_1431_io_cout; // @[MUL.scala 253:22]
  assign m_1773_io_x3 = m_1436_io_s; // @[MUL.scala 252:21]
  assign m_1774_io_x1 = m_1432_io_cout; // @[MUL.scala 253:22]
  assign m_1774_io_x2 = m_1437_io_s; // @[MUL.scala 252:21]
  assign m_1774_io_x3 = m_1433_io_cout; // @[MUL.scala 253:22]
  assign m_1775_io_in_0 = m_1438_io_s; // @[MUL.scala 252:21]
  assign m_1775_io_in_1 = m_1434_io_cout; // @[MUL.scala 253:22]
  assign m_1776_io_x1 = m_1439_io_s; // @[MUL.scala 252:21]
  assign m_1776_io_x2 = m_1435_io_cout; // @[MUL.scala 253:22]
  assign m_1776_io_x3 = m_1440_io_s; // @[MUL.scala 252:21]
  assign m_1777_io_x1 = m_1436_io_cout; // @[MUL.scala 253:22]
  assign m_1777_io_x2 = m_1441_io_s; // @[MUL.scala 252:21]
  assign m_1777_io_x3 = m_1437_io_cout; // @[MUL.scala 253:22]
  assign m_1778_io_in_0 = m_1442_io_s; // @[MUL.scala 252:21]
  assign m_1778_io_in_1 = m_1438_io_cout; // @[MUL.scala 253:22]
  assign m_1779_io_x1 = m_1443_io_s; // @[MUL.scala 252:21]
  assign m_1779_io_x2 = m_1439_io_cout; // @[MUL.scala 253:22]
  assign m_1779_io_x3 = m_1444_io_s; // @[MUL.scala 252:21]
  assign m_1780_io_x1 = m_1440_io_cout; // @[MUL.scala 253:22]
  assign m_1780_io_x2 = m_1445_io_s; // @[MUL.scala 252:21]
  assign m_1780_io_x3 = m_1441_io_cout; // @[MUL.scala 253:22]
  assign m_1781_io_in_0 = m_1446_io_s; // @[MUL.scala 252:21]
  assign m_1781_io_in_1 = m_1442_io_cout; // @[MUL.scala 253:22]
  assign m_1782_io_x1 = m_1447_io_s; // @[MUL.scala 252:21]
  assign m_1782_io_x2 = m_1443_io_cout; // @[MUL.scala 253:22]
  assign m_1782_io_x3 = m_1448_io_s; // @[MUL.scala 252:21]
  assign m_1783_io_x1 = m_1444_io_cout; // @[MUL.scala 253:22]
  assign m_1783_io_x2 = m_1449_io_s; // @[MUL.scala 252:21]
  assign m_1783_io_x3 = m_1445_io_cout; // @[MUL.scala 253:22]
  assign m_1784_io_x1 = m_1450_io_s; // @[MUL.scala 252:21]
  assign m_1784_io_x2 = m_1446_io_cout; // @[MUL.scala 253:22]
  assign m_1784_io_x3 = r_781; // @[MUL.scala 105:13]
  assign m_1785_io_x1 = m_1451_io_s; // @[MUL.scala 252:21]
  assign m_1785_io_x2 = m_1447_io_cout; // @[MUL.scala 253:22]
  assign m_1785_io_x3 = m_1452_io_s; // @[MUL.scala 252:21]
  assign m_1786_io_x1 = m_1448_io_cout; // @[MUL.scala 253:22]
  assign m_1786_io_x2 = m_1453_io_s; // @[MUL.scala 252:21]
  assign m_1786_io_x3 = m_1449_io_cout; // @[MUL.scala 253:22]
  assign m_1787_io_x1 = m_1454_io_s; // @[MUL.scala 252:21]
  assign m_1787_io_x2 = m_1450_io_cout; // @[MUL.scala 253:22]
  assign m_1787_io_x3 = r_809; // @[MUL.scala 105:13]
  assign m_1788_io_x1 = m_1455_io_s; // @[MUL.scala 252:21]
  assign m_1788_io_x2 = m_1451_io_cout; // @[MUL.scala 253:22]
  assign m_1788_io_x3 = m_1456_io_s; // @[MUL.scala 252:21]
  assign m_1789_io_x1 = m_1452_io_cout; // @[MUL.scala 253:22]
  assign m_1789_io_x2 = m_1457_io_s; // @[MUL.scala 252:21]
  assign m_1789_io_x3 = m_1453_io_cout; // @[MUL.scala 253:22]
  assign m_1790_io_x1 = m_1458_io_s; // @[MUL.scala 252:21]
  assign m_1790_io_x2 = m_1454_io_cout; // @[MUL.scala 253:22]
  assign m_1790_io_x3 = m_312_io_out_0; // @[MUL.scala 105:13]
  assign m_1791_io_x1 = m_1459_io_s; // @[MUL.scala 252:21]
  assign m_1791_io_x2 = m_1455_io_cout; // @[MUL.scala 253:22]
  assign m_1791_io_x3 = m_1460_io_s; // @[MUL.scala 252:21]
  assign m_1792_io_x1 = m_1456_io_cout; // @[MUL.scala 253:22]
  assign m_1792_io_x2 = m_1461_io_s; // @[MUL.scala 252:21]
  assign m_1792_io_x3 = m_1457_io_cout; // @[MUL.scala 253:22]
  assign m_1793_io_x1 = m_1462_io_s; // @[MUL.scala 252:21]
  assign m_1793_io_x2 = m_1458_io_cout; // @[MUL.scala 253:22]
  assign m_1793_io_x3 = m_998_io_out_0; // @[MUL.scala 105:13]
  assign m_1794_io_x1 = m_1463_io_s; // @[MUL.scala 252:21]
  assign m_1794_io_x2 = m_1459_io_cout; // @[MUL.scala 253:22]
  assign m_1794_io_x3 = m_1464_io_s; // @[MUL.scala 252:21]
  assign m_1795_io_x1 = m_1460_io_cout; // @[MUL.scala 253:22]
  assign m_1795_io_x2 = m_1465_io_s; // @[MUL.scala 252:21]
  assign m_1795_io_x3 = m_1461_io_cout; // @[MUL.scala 253:22]
  assign m_1796_io_x1 = m_1466_io_s; // @[MUL.scala 252:21]
  assign m_1796_io_x2 = m_1462_io_cout; // @[MUL.scala 253:22]
  assign m_1796_io_x3 = m_1467_io_out_0; // @[MUL.scala 105:13]
  assign m_1797_io_x1 = m_1468_io_s; // @[MUL.scala 252:21]
  assign m_1797_io_x2 = m_1463_io_cout; // @[MUL.scala 253:22]
  assign m_1797_io_x3 = m_1469_io_s; // @[MUL.scala 252:21]
  assign m_1798_io_x1 = m_1464_io_cout; // @[MUL.scala 253:22]
  assign m_1798_io_x2 = m_1470_io_s; // @[MUL.scala 252:21]
  assign m_1798_io_x3 = m_1465_io_cout; // @[MUL.scala 253:22]
  assign m_1799_io_x1 = m_1471_io_s; // @[MUL.scala 252:21]
  assign m_1799_io_x2 = m_1466_io_cout; // @[MUL.scala 253:22]
  assign m_1799_io_x3 = m_1472_io_out_0; // @[MUL.scala 105:13]
  assign m_1800_io_x1 = m_1473_io_s; // @[MUL.scala 252:21]
  assign m_1800_io_x2 = m_1468_io_cout; // @[MUL.scala 253:22]
  assign m_1800_io_x3 = m_1474_io_s; // @[MUL.scala 252:21]
  assign m_1801_io_x1 = m_1469_io_cout; // @[MUL.scala 253:22]
  assign m_1801_io_x2 = m_1475_io_s; // @[MUL.scala 252:21]
  assign m_1801_io_x3 = m_1470_io_cout; // @[MUL.scala 253:22]
  assign m_1802_io_x1 = m_1476_io_s; // @[MUL.scala 252:21]
  assign m_1802_io_x2 = m_1471_io_cout; // @[MUL.scala 253:22]
  assign m_1802_io_x3 = m_1477_io_out_0; // @[MUL.scala 105:13]
  assign m_1803_io_x1 = m_1478_io_s; // @[MUL.scala 252:21]
  assign m_1803_io_x2 = m_1473_io_cout; // @[MUL.scala 253:22]
  assign m_1803_io_x3 = m_1479_io_s; // @[MUL.scala 252:21]
  assign m_1804_io_x1 = m_1474_io_cout; // @[MUL.scala 253:22]
  assign m_1804_io_x2 = m_1480_io_s; // @[MUL.scala 252:21]
  assign m_1804_io_x3 = m_1475_io_cout; // @[MUL.scala 253:22]
  assign m_1805_io_x1 = m_1481_io_s; // @[MUL.scala 252:21]
  assign m_1805_io_x2 = m_1476_io_cout; // @[MUL.scala 253:22]
  assign m_1805_io_x3 = m_1482_io_out_0; // @[MUL.scala 105:13]
  assign m_1806_io_x1 = m_1483_io_s; // @[MUL.scala 252:21]
  assign m_1806_io_x2 = m_1478_io_cout; // @[MUL.scala 253:22]
  assign m_1806_io_x3 = m_1484_io_s; // @[MUL.scala 252:21]
  assign m_1807_io_x1 = m_1479_io_cout; // @[MUL.scala 253:22]
  assign m_1807_io_x2 = m_1485_io_s; // @[MUL.scala 252:21]
  assign m_1807_io_x3 = m_1480_io_cout; // @[MUL.scala 253:22]
  assign m_1808_io_x1 = m_1486_io_s; // @[MUL.scala 252:21]
  assign m_1808_io_x2 = m_1481_io_cout; // @[MUL.scala 253:22]
  assign m_1808_io_x3 = m_1487_io_out_0; // @[MUL.scala 105:13]
  assign m_1809_io_x1 = m_1488_io_s; // @[MUL.scala 252:21]
  assign m_1809_io_x2 = m_1483_io_cout; // @[MUL.scala 253:22]
  assign m_1809_io_x3 = m_1489_io_s; // @[MUL.scala 252:21]
  assign m_1810_io_x1 = m_1484_io_cout; // @[MUL.scala 253:22]
  assign m_1810_io_x2 = m_1490_io_s; // @[MUL.scala 252:21]
  assign m_1810_io_x3 = m_1485_io_cout; // @[MUL.scala 253:22]
  assign m_1811_io_x1 = m_1491_io_s; // @[MUL.scala 252:21]
  assign m_1811_io_x2 = m_1486_io_cout; // @[MUL.scala 253:22]
  assign m_1811_io_x3 = m_1492_io_s; // @[MUL.scala 252:21]
  assign m_1812_io_x1 = m_1493_io_s; // @[MUL.scala 252:21]
  assign m_1812_io_x2 = m_1488_io_cout; // @[MUL.scala 253:22]
  assign m_1812_io_x3 = m_1494_io_s; // @[MUL.scala 252:21]
  assign m_1813_io_x1 = m_1489_io_cout; // @[MUL.scala 253:22]
  assign m_1813_io_x2 = m_1495_io_s; // @[MUL.scala 252:21]
  assign m_1813_io_x3 = m_1490_io_cout; // @[MUL.scala 253:22]
  assign m_1814_io_x1 = m_1496_io_s; // @[MUL.scala 252:21]
  assign m_1814_io_x2 = m_1491_io_cout; // @[MUL.scala 253:22]
  assign m_1814_io_x3 = m_1497_io_s; // @[MUL.scala 252:21]
  assign m_1815_io_x1 = m_1498_io_s; // @[MUL.scala 252:21]
  assign m_1815_io_x2 = m_1493_io_cout; // @[MUL.scala 253:22]
  assign m_1815_io_x3 = m_1499_io_s; // @[MUL.scala 252:21]
  assign m_1816_io_x1 = m_1494_io_cout; // @[MUL.scala 253:22]
  assign m_1816_io_x2 = m_1500_io_s; // @[MUL.scala 252:21]
  assign m_1816_io_x3 = m_1495_io_cout; // @[MUL.scala 253:22]
  assign m_1817_io_x1 = m_1501_io_s; // @[MUL.scala 252:21]
  assign m_1817_io_x2 = m_1496_io_cout; // @[MUL.scala 253:22]
  assign m_1817_io_x3 = m_1502_io_s; // @[MUL.scala 252:21]
  assign m_1818_io_x1 = m_1503_io_s; // @[MUL.scala 252:21]
  assign m_1818_io_x2 = m_1498_io_cout; // @[MUL.scala 253:22]
  assign m_1818_io_x3 = m_1504_io_s; // @[MUL.scala 252:21]
  assign m_1819_io_x1 = m_1499_io_cout; // @[MUL.scala 253:22]
  assign m_1819_io_x2 = m_1505_io_s; // @[MUL.scala 252:21]
  assign m_1819_io_x3 = m_1500_io_cout; // @[MUL.scala 253:22]
  assign m_1820_io_x1 = m_1506_io_s; // @[MUL.scala 252:21]
  assign m_1820_io_x2 = m_1501_io_cout; // @[MUL.scala 253:22]
  assign m_1820_io_x3 = m_1507_io_s; // @[MUL.scala 252:21]
  assign m_1821_io_x1 = m_1508_io_s; // @[MUL.scala 252:21]
  assign m_1821_io_x2 = m_1503_io_cout; // @[MUL.scala 253:22]
  assign m_1821_io_x3 = m_1509_io_s; // @[MUL.scala 252:21]
  assign m_1822_io_x1 = m_1504_io_cout; // @[MUL.scala 253:22]
  assign m_1822_io_x2 = m_1510_io_s; // @[MUL.scala 252:21]
  assign m_1822_io_x3 = m_1505_io_cout; // @[MUL.scala 253:22]
  assign m_1823_io_x1 = m_1511_io_s; // @[MUL.scala 252:21]
  assign m_1823_io_x2 = m_1506_io_cout; // @[MUL.scala 253:22]
  assign m_1823_io_x3 = m_1512_io_s; // @[MUL.scala 252:21]
  assign m_1824_io_x1 = m_1513_io_s; // @[MUL.scala 252:21]
  assign m_1824_io_x2 = m_1508_io_cout; // @[MUL.scala 253:22]
  assign m_1824_io_x3 = m_1514_io_s; // @[MUL.scala 252:21]
  assign m_1825_io_x1 = m_1509_io_cout; // @[MUL.scala 253:22]
  assign m_1825_io_x2 = m_1515_io_s; // @[MUL.scala 252:21]
  assign m_1825_io_x3 = m_1510_io_cout; // @[MUL.scala 253:22]
  assign m_1826_io_x1 = m_1516_io_s; // @[MUL.scala 252:21]
  assign m_1826_io_x2 = m_1511_io_cout; // @[MUL.scala 253:22]
  assign m_1826_io_x3 = m_1517_io_s; // @[MUL.scala 252:21]
  assign m_1827_io_x1 = m_1518_io_s; // @[MUL.scala 252:21]
  assign m_1827_io_x2 = m_1513_io_cout; // @[MUL.scala 253:22]
  assign m_1827_io_x3 = m_1519_io_s; // @[MUL.scala 252:21]
  assign m_1828_io_x1 = m_1514_io_cout; // @[MUL.scala 253:22]
  assign m_1828_io_x2 = m_1520_io_s; // @[MUL.scala 252:21]
  assign m_1828_io_x3 = m_1515_io_cout; // @[MUL.scala 253:22]
  assign m_1829_io_x1 = m_1521_io_s; // @[MUL.scala 252:21]
  assign m_1829_io_x2 = m_1516_io_cout; // @[MUL.scala 253:22]
  assign m_1829_io_x3 = m_1522_io_s; // @[MUL.scala 252:21]
  assign m_1830_io_x1 = m_1523_io_s; // @[MUL.scala 252:21]
  assign m_1830_io_x2 = m_1518_io_cout; // @[MUL.scala 253:22]
  assign m_1830_io_x3 = m_1524_io_s; // @[MUL.scala 252:21]
  assign m_1831_io_x1 = m_1519_io_cout; // @[MUL.scala 253:22]
  assign m_1831_io_x2 = m_1525_io_s; // @[MUL.scala 252:21]
  assign m_1831_io_x3 = m_1520_io_cout; // @[MUL.scala 253:22]
  assign m_1832_io_x1 = m_1526_io_s; // @[MUL.scala 252:21]
  assign m_1832_io_x2 = m_1521_io_cout; // @[MUL.scala 253:22]
  assign m_1832_io_x3 = m_1527_io_s; // @[MUL.scala 252:21]
  assign m_1833_io_x1 = m_1528_io_s; // @[MUL.scala 252:21]
  assign m_1833_io_x2 = m_1523_io_cout; // @[MUL.scala 253:22]
  assign m_1833_io_x3 = m_1529_io_s; // @[MUL.scala 252:21]
  assign m_1834_io_x1 = m_1524_io_cout; // @[MUL.scala 253:22]
  assign m_1834_io_x2 = m_1530_io_s; // @[MUL.scala 252:21]
  assign m_1834_io_x3 = m_1525_io_cout; // @[MUL.scala 253:22]
  assign m_1835_io_x1 = m_1531_io_s; // @[MUL.scala 252:21]
  assign m_1835_io_x2 = m_1526_io_cout; // @[MUL.scala 253:22]
  assign m_1835_io_x3 = m_1532_io_s; // @[MUL.scala 252:21]
  assign m_1836_io_x1 = m_1533_io_s; // @[MUL.scala 252:21]
  assign m_1836_io_x2 = m_1528_io_cout; // @[MUL.scala 253:22]
  assign m_1836_io_x3 = m_1534_io_s; // @[MUL.scala 252:21]
  assign m_1837_io_x1 = m_1529_io_cout; // @[MUL.scala 253:22]
  assign m_1837_io_x2 = m_1535_io_s; // @[MUL.scala 252:21]
  assign m_1837_io_x3 = m_1530_io_cout; // @[MUL.scala 253:22]
  assign m_1838_io_x1 = m_1536_io_s; // @[MUL.scala 252:21]
  assign m_1838_io_x2 = m_1531_io_cout; // @[MUL.scala 253:22]
  assign m_1838_io_x3 = m_1537_io_s; // @[MUL.scala 252:21]
  assign m_1839_io_x1 = m_1538_io_s; // @[MUL.scala 252:21]
  assign m_1839_io_x2 = m_1533_io_cout; // @[MUL.scala 253:22]
  assign m_1839_io_x3 = m_1539_io_s; // @[MUL.scala 252:21]
  assign m_1840_io_x1 = m_1534_io_cout; // @[MUL.scala 253:22]
  assign m_1840_io_x2 = m_1540_io_s; // @[MUL.scala 252:21]
  assign m_1840_io_x3 = m_1535_io_cout; // @[MUL.scala 253:22]
  assign m_1841_io_x1 = m_1541_io_s; // @[MUL.scala 252:21]
  assign m_1841_io_x2 = m_1536_io_cout; // @[MUL.scala 253:22]
  assign m_1841_io_x3 = m_1542_io_out_0; // @[MUL.scala 105:13]
  assign m_1842_io_x1 = m_1543_io_s; // @[MUL.scala 252:21]
  assign m_1842_io_x2 = m_1538_io_cout; // @[MUL.scala 253:22]
  assign m_1842_io_x3 = m_1544_io_s; // @[MUL.scala 252:21]
  assign m_1843_io_x1 = m_1539_io_cout; // @[MUL.scala 253:22]
  assign m_1843_io_x2 = m_1545_io_s; // @[MUL.scala 252:21]
  assign m_1843_io_x3 = m_1540_io_cout; // @[MUL.scala 253:22]
  assign m_1844_io_x1 = m_1546_io_s; // @[MUL.scala 252:21]
  assign m_1844_io_x2 = m_1541_io_cout; // @[MUL.scala 253:22]
  assign m_1844_io_x3 = m_1547_io_out_0; // @[MUL.scala 105:13]
  assign m_1845_io_x1 = m_1548_io_s; // @[MUL.scala 252:21]
  assign m_1845_io_x2 = m_1543_io_cout; // @[MUL.scala 253:22]
  assign m_1845_io_x3 = m_1549_io_s; // @[MUL.scala 252:21]
  assign m_1846_io_x1 = m_1544_io_cout; // @[MUL.scala 253:22]
  assign m_1846_io_x2 = m_1550_io_s; // @[MUL.scala 252:21]
  assign m_1846_io_x3 = m_1545_io_cout; // @[MUL.scala 253:22]
  assign m_1847_io_x1 = m_1551_io_s; // @[MUL.scala 252:21]
  assign m_1847_io_x2 = m_1546_io_cout; // @[MUL.scala 253:22]
  assign m_1847_io_x3 = m_1552_io_out_0; // @[MUL.scala 105:13]
  assign m_1848_io_x1 = m_1553_io_s; // @[MUL.scala 252:21]
  assign m_1848_io_x2 = m_1548_io_cout; // @[MUL.scala 253:22]
  assign m_1848_io_x3 = m_1554_io_s; // @[MUL.scala 252:21]
  assign m_1849_io_x1 = m_1549_io_cout; // @[MUL.scala 253:22]
  assign m_1849_io_x2 = m_1555_io_s; // @[MUL.scala 252:21]
  assign m_1849_io_x3 = m_1550_io_cout; // @[MUL.scala 253:22]
  assign m_1850_io_x1 = m_1556_io_s; // @[MUL.scala 252:21]
  assign m_1850_io_x2 = m_1551_io_cout; // @[MUL.scala 253:22]
  assign m_1850_io_x3 = m_1557_io_out_0; // @[MUL.scala 105:13]
  assign m_1851_io_x1 = m_1558_io_s; // @[MUL.scala 252:21]
  assign m_1851_io_x2 = m_1553_io_cout; // @[MUL.scala 253:22]
  assign m_1851_io_x3 = m_1559_io_s; // @[MUL.scala 252:21]
  assign m_1852_io_x1 = m_1554_io_cout; // @[MUL.scala 253:22]
  assign m_1852_io_x2 = m_1560_io_s; // @[MUL.scala 252:21]
  assign m_1852_io_x3 = m_1555_io_cout; // @[MUL.scala 253:22]
  assign m_1853_io_x1 = m_1561_io_s; // @[MUL.scala 252:21]
  assign m_1853_io_x2 = m_1556_io_cout; // @[MUL.scala 253:22]
  assign m_1853_io_x3 = m_1562_io_out_0; // @[MUL.scala 105:13]
  assign m_1854_io_x1 = m_1563_io_s; // @[MUL.scala 252:21]
  assign m_1854_io_x2 = m_1558_io_cout; // @[MUL.scala 253:22]
  assign m_1854_io_x3 = m_1564_io_s; // @[MUL.scala 252:21]
  assign m_1855_io_x1 = m_1559_io_cout; // @[MUL.scala 253:22]
  assign m_1855_io_x2 = m_1565_io_s; // @[MUL.scala 252:21]
  assign m_1855_io_x3 = m_1560_io_cout; // @[MUL.scala 253:22]
  assign m_1856_io_x1 = m_1566_io_s; // @[MUL.scala 252:21]
  assign m_1856_io_x2 = m_1561_io_cout; // @[MUL.scala 253:22]
  assign m_1856_io_x3 = m_1567_io_out_0; // @[MUL.scala 105:13]
  assign m_1857_io_x1 = m_1568_io_s; // @[MUL.scala 252:21]
  assign m_1857_io_x2 = m_1563_io_cout; // @[MUL.scala 253:22]
  assign m_1857_io_x3 = m_1569_io_s; // @[MUL.scala 252:21]
  assign m_1858_io_x1 = m_1564_io_cout; // @[MUL.scala 253:22]
  assign m_1858_io_x2 = m_1570_io_s; // @[MUL.scala 252:21]
  assign m_1858_io_x3 = m_1565_io_cout; // @[MUL.scala 253:22]
  assign m_1859_io_x1 = m_1571_io_s; // @[MUL.scala 252:21]
  assign m_1859_io_x2 = m_1566_io_cout; // @[MUL.scala 253:22]
  assign m_1859_io_x3 = m_1572_io_out_0; // @[MUL.scala 105:13]
  assign m_1860_io_x1 = m_1573_io_s; // @[MUL.scala 252:21]
  assign m_1860_io_x2 = m_1568_io_cout; // @[MUL.scala 253:22]
  assign m_1860_io_x3 = m_1574_io_s; // @[MUL.scala 252:21]
  assign m_1861_io_x1 = m_1569_io_cout; // @[MUL.scala 253:22]
  assign m_1861_io_x2 = m_1575_io_s; // @[MUL.scala 252:21]
  assign m_1861_io_x3 = m_1570_io_cout; // @[MUL.scala 253:22]
  assign m_1862_io_x1 = m_1576_io_s; // @[MUL.scala 252:21]
  assign m_1862_io_x2 = m_1571_io_cout; // @[MUL.scala 253:22]
  assign m_1862_io_x3 = m_1572_io_out_1; // @[MUL.scala 105:13]
  assign m_1863_io_x1 = m_1577_io_s; // @[MUL.scala 252:21]
  assign m_1863_io_x2 = m_1573_io_cout; // @[MUL.scala 253:22]
  assign m_1863_io_x3 = m_1578_io_s; // @[MUL.scala 252:21]
  assign m_1864_io_x1 = m_1574_io_cout; // @[MUL.scala 253:22]
  assign m_1864_io_x2 = m_1579_io_s; // @[MUL.scala 252:21]
  assign m_1864_io_x3 = m_1575_io_cout; // @[MUL.scala 253:22]
  assign m_1865_io_in_0 = m_1580_io_s; // @[MUL.scala 252:21]
  assign m_1865_io_in_1 = m_1576_io_cout; // @[MUL.scala 253:22]
  assign m_1866_io_x1 = m_1581_io_s; // @[MUL.scala 252:21]
  assign m_1866_io_x2 = m_1577_io_cout; // @[MUL.scala 253:22]
  assign m_1866_io_x3 = m_1582_io_s; // @[MUL.scala 252:21]
  assign m_1867_io_x1 = m_1578_io_cout; // @[MUL.scala 253:22]
  assign m_1867_io_x2 = m_1583_io_s; // @[MUL.scala 252:21]
  assign m_1867_io_x3 = m_1579_io_cout; // @[MUL.scala 253:22]
  assign m_1868_io_in_0 = m_1584_io_s; // @[MUL.scala 252:21]
  assign m_1868_io_in_1 = m_1580_io_cout; // @[MUL.scala 253:22]
  assign m_1869_io_x1 = m_1585_io_s; // @[MUL.scala 252:21]
  assign m_1869_io_x2 = m_1581_io_cout; // @[MUL.scala 253:22]
  assign m_1869_io_x3 = m_1586_io_s; // @[MUL.scala 252:21]
  assign m_1870_io_x1 = m_1582_io_cout; // @[MUL.scala 253:22]
  assign m_1870_io_x2 = m_1587_io_s; // @[MUL.scala 252:21]
  assign m_1870_io_x3 = m_1583_io_cout; // @[MUL.scala 253:22]
  assign m_1871_io_in_0 = m_1588_io_s; // @[MUL.scala 252:21]
  assign m_1871_io_in_1 = m_1584_io_cout; // @[MUL.scala 253:22]
  assign m_1872_io_x1 = m_1589_io_s; // @[MUL.scala 252:21]
  assign m_1872_io_x2 = m_1585_io_cout; // @[MUL.scala 253:22]
  assign m_1872_io_x3 = m_1590_io_s; // @[MUL.scala 252:21]
  assign m_1873_io_x1 = m_1586_io_cout; // @[MUL.scala 253:22]
  assign m_1873_io_x2 = m_1591_io_s; // @[MUL.scala 252:21]
  assign m_1873_io_x3 = m_1587_io_cout; // @[MUL.scala 253:22]
  assign m_1874_io_in_0 = m_1592_io_s; // @[MUL.scala 252:21]
  assign m_1874_io_in_1 = m_1588_io_cout; // @[MUL.scala 253:22]
  assign m_1875_io_x1 = m_1593_io_s; // @[MUL.scala 252:21]
  assign m_1875_io_x2 = m_1589_io_cout; // @[MUL.scala 253:22]
  assign m_1875_io_x3 = m_1594_io_s; // @[MUL.scala 252:21]
  assign m_1876_io_x1 = m_1590_io_cout; // @[MUL.scala 253:22]
  assign m_1876_io_x2 = m_1595_io_s; // @[MUL.scala 252:21]
  assign m_1876_io_x3 = m_1591_io_cout; // @[MUL.scala 253:22]
  assign m_1877_io_in_0 = m_1596_io_s; // @[MUL.scala 252:21]
  assign m_1877_io_in_1 = m_1592_io_cout; // @[MUL.scala 253:22]
  assign m_1878_io_x1 = m_1597_io_s; // @[MUL.scala 252:21]
  assign m_1878_io_x2 = m_1593_io_cout; // @[MUL.scala 253:22]
  assign m_1878_io_x3 = m_1598_io_s; // @[MUL.scala 252:21]
  assign m_1879_io_x1 = m_1594_io_cout; // @[MUL.scala 253:22]
  assign m_1879_io_x2 = m_1599_io_s; // @[MUL.scala 252:21]
  assign m_1879_io_x3 = m_1595_io_cout; // @[MUL.scala 253:22]
  assign m_1880_io_in_0 = m_1600_io_s; // @[MUL.scala 252:21]
  assign m_1880_io_in_1 = m_1596_io_cout; // @[MUL.scala 253:22]
  assign m_1881_io_x1 = m_1601_io_s; // @[MUL.scala 252:21]
  assign m_1881_io_x2 = m_1597_io_cout; // @[MUL.scala 253:22]
  assign m_1881_io_x3 = m_1602_io_s; // @[MUL.scala 252:21]
  assign m_1882_io_x1 = m_1598_io_cout; // @[MUL.scala 253:22]
  assign m_1882_io_x2 = m_1603_io_s; // @[MUL.scala 252:21]
  assign m_1882_io_x3 = m_1599_io_cout; // @[MUL.scala 253:22]
  assign m_1883_io_in_0 = m_1604_io_out_0; // @[MUL.scala 125:16]
  assign m_1883_io_in_1 = m_1600_io_cout; // @[MUL.scala 253:22]
  assign m_1884_io_x1 = m_1605_io_s; // @[MUL.scala 252:21]
  assign m_1884_io_x2 = m_1601_io_cout; // @[MUL.scala 253:22]
  assign m_1884_io_x3 = m_1606_io_s; // @[MUL.scala 252:21]
  assign m_1885_io_x1 = m_1602_io_cout; // @[MUL.scala 253:22]
  assign m_1885_io_x2 = m_1607_io_s; // @[MUL.scala 252:21]
  assign m_1885_io_x3 = m_1603_io_cout; // @[MUL.scala 253:22]
  assign m_1886_io_in_0 = m_1608_io_out_0; // @[MUL.scala 125:16]
  assign m_1886_io_in_1 = m_1604_io_out_1; // @[MUL.scala 126:16]
  assign m_1887_io_x1 = m_1609_io_s; // @[MUL.scala 252:21]
  assign m_1887_io_x2 = m_1605_io_cout; // @[MUL.scala 253:22]
  assign m_1887_io_x3 = m_1610_io_s; // @[MUL.scala 252:21]
  assign m_1888_io_x1 = m_1606_io_cout; // @[MUL.scala 253:22]
  assign m_1888_io_x2 = m_1611_io_s; // @[MUL.scala 252:21]
  assign m_1888_io_x3 = m_1607_io_cout; // @[MUL.scala 253:22]
  assign m_1889_io_in_0 = m_1612_io_out_0; // @[MUL.scala 125:16]
  assign m_1889_io_in_1 = m_1608_io_out_1; // @[MUL.scala 126:16]
  assign m_1890_io_x1 = m_1613_io_s; // @[MUL.scala 252:21]
  assign m_1890_io_x2 = m_1609_io_cout; // @[MUL.scala 253:22]
  assign m_1890_io_x3 = m_1614_io_s; // @[MUL.scala 252:21]
  assign m_1891_io_x1 = m_1610_io_cout; // @[MUL.scala 253:22]
  assign m_1891_io_x2 = m_1615_io_s; // @[MUL.scala 252:21]
  assign m_1891_io_x3 = m_1611_io_cout; // @[MUL.scala 253:22]
  assign m_1892_io_in_0 = m_1616_io_out_0; // @[MUL.scala 125:16]
  assign m_1892_io_in_1 = m_1612_io_out_1; // @[MUL.scala 126:16]
  assign m_1893_io_x1 = m_1617_io_s; // @[MUL.scala 252:21]
  assign m_1893_io_x2 = m_1613_io_cout; // @[MUL.scala 253:22]
  assign m_1893_io_x3 = m_1618_io_s; // @[MUL.scala 252:21]
  assign m_1894_io_x1 = m_1614_io_cout; // @[MUL.scala 253:22]
  assign m_1894_io_x2 = m_1619_io_s; // @[MUL.scala 252:21]
  assign m_1894_io_x3 = m_1615_io_cout; // @[MUL.scala 253:22]
  assign m_1895_io_in_0 = m_1212_io_cout; // @[MUL.scala 253:22]
  assign m_1895_io_in_1 = m_1616_io_out_1; // @[MUL.scala 126:16]
  assign m_1896_io_x1 = m_1620_io_s; // @[MUL.scala 252:21]
  assign m_1896_io_x2 = m_1617_io_cout; // @[MUL.scala 253:22]
  assign m_1896_io_x3 = m_1621_io_s; // @[MUL.scala 252:21]
  assign m_1897_io_x1 = m_1618_io_cout; // @[MUL.scala 253:22]
  assign m_1897_io_x2 = m_1622_io_s; // @[MUL.scala 252:21]
  assign m_1897_io_x3 = m_1619_io_cout; // @[MUL.scala 253:22]
  assign m_1898_io_x1 = m_1623_io_s; // @[MUL.scala 252:21]
  assign m_1898_io_x2 = m_1620_io_cout; // @[MUL.scala 253:22]
  assign m_1898_io_x3 = m_1624_io_s; // @[MUL.scala 252:21]
  assign m_1899_io_x1 = m_1621_io_cout; // @[MUL.scala 253:22]
  assign m_1899_io_x2 = m_1625_io_s; // @[MUL.scala 252:21]
  assign m_1899_io_x3 = m_1622_io_cout; // @[MUL.scala 253:22]
  assign m_1900_io_x1 = m_1626_io_s; // @[MUL.scala 252:21]
  assign m_1900_io_x2 = m_1623_io_cout; // @[MUL.scala 253:22]
  assign m_1900_io_x3 = m_1627_io_s; // @[MUL.scala 252:21]
  assign m_1901_io_x1 = m_1624_io_cout; // @[MUL.scala 253:22]
  assign m_1901_io_x2 = m_1628_io_s; // @[MUL.scala 252:21]
  assign m_1901_io_x3 = m_1625_io_cout; // @[MUL.scala 253:22]
  assign m_1902_io_x1 = m_1629_io_s; // @[MUL.scala 252:21]
  assign m_1902_io_x2 = m_1626_io_cout; // @[MUL.scala 253:22]
  assign m_1902_io_x3 = m_1630_io_s; // @[MUL.scala 252:21]
  assign m_1903_io_x1 = m_1627_io_cout; // @[MUL.scala 253:22]
  assign m_1903_io_x2 = m_1631_io_s; // @[MUL.scala 252:21]
  assign m_1903_io_x3 = m_1628_io_cout; // @[MUL.scala 253:22]
  assign m_1904_io_x1 = m_1632_io_s; // @[MUL.scala 252:21]
  assign m_1904_io_x2 = m_1629_io_cout; // @[MUL.scala 253:22]
  assign m_1904_io_x3 = m_1633_io_s; // @[MUL.scala 252:21]
  assign m_1905_io_x1 = m_1630_io_cout; // @[MUL.scala 253:22]
  assign m_1905_io_x2 = m_1634_io_s; // @[MUL.scala 252:21]
  assign m_1905_io_x3 = m_1631_io_cout; // @[MUL.scala 253:22]
  assign m_1906_io_x1 = m_1635_io_s; // @[MUL.scala 252:21]
  assign m_1906_io_x2 = m_1632_io_cout; // @[MUL.scala 253:22]
  assign m_1906_io_x3 = m_1636_io_s; // @[MUL.scala 252:21]
  assign m_1907_io_x1 = m_1633_io_cout; // @[MUL.scala 253:22]
  assign m_1907_io_x2 = m_1637_io_s; // @[MUL.scala 252:21]
  assign m_1907_io_x3 = m_1634_io_cout; // @[MUL.scala 253:22]
  assign m_1908_io_x1 = m_1638_io_s; // @[MUL.scala 252:21]
  assign m_1908_io_x2 = m_1635_io_cout; // @[MUL.scala 253:22]
  assign m_1908_io_x3 = m_1639_io_s; // @[MUL.scala 252:21]
  assign m_1909_io_x1 = m_1636_io_cout; // @[MUL.scala 253:22]
  assign m_1909_io_x2 = m_1640_io_out_0; // @[MUL.scala 104:13]
  assign m_1909_io_x3 = m_1637_io_cout; // @[MUL.scala 253:22]
  assign m_1910_io_x1 = m_1641_io_s; // @[MUL.scala 252:21]
  assign m_1910_io_x2 = m_1638_io_cout; // @[MUL.scala 253:22]
  assign m_1910_io_x3 = m_1642_io_s; // @[MUL.scala 252:21]
  assign m_1911_io_x1 = m_1639_io_cout; // @[MUL.scala 253:22]
  assign m_1911_io_x2 = m_1643_io_out_0; // @[MUL.scala 104:13]
  assign m_1911_io_x3 = m_1640_io_out_1; // @[MUL.scala 105:13]
  assign m_1912_io_x1 = m_1644_io_s; // @[MUL.scala 252:21]
  assign m_1912_io_x2 = m_1641_io_cout; // @[MUL.scala 253:22]
  assign m_1912_io_x3 = m_1645_io_s; // @[MUL.scala 252:21]
  assign m_1913_io_x1 = m_1642_io_cout; // @[MUL.scala 253:22]
  assign m_1913_io_x2 = m_1646_io_out_0; // @[MUL.scala 104:13]
  assign m_1913_io_x3 = m_1643_io_out_1; // @[MUL.scala 105:13]
  assign m_1914_io_x1 = m_1647_io_s; // @[MUL.scala 252:21]
  assign m_1914_io_x2 = m_1644_io_cout; // @[MUL.scala 253:22]
  assign m_1914_io_x3 = m_1648_io_s; // @[MUL.scala 252:21]
  assign m_1915_io_x1 = m_1645_io_cout; // @[MUL.scala 253:22]
  assign m_1915_io_x2 = m_1649_io_out_0; // @[MUL.scala 104:13]
  assign m_1915_io_x3 = m_1646_io_out_1; // @[MUL.scala 105:13]
  assign m_1916_io_x1 = m_1650_io_s; // @[MUL.scala 252:21]
  assign m_1916_io_x2 = m_1647_io_cout; // @[MUL.scala 253:22]
  assign m_1916_io_x3 = m_1651_io_s; // @[MUL.scala 252:21]
  assign m_1917_io_x1 = m_1648_io_cout; // @[MUL.scala 253:22]
  assign m_1917_io_x2 = m_1652_io_out_0; // @[MUL.scala 104:13]
  assign m_1917_io_x3 = m_1649_io_out_1; // @[MUL.scala 105:13]
  assign m_1918_io_x1 = m_1653_io_s; // @[MUL.scala 252:21]
  assign m_1918_io_x2 = m_1650_io_cout; // @[MUL.scala 253:22]
  assign m_1918_io_x3 = m_1654_io_s; // @[MUL.scala 252:21]
  assign m_1919_io_x1 = m_1651_io_cout; // @[MUL.scala 253:22]
  assign m_1919_io_x2 = m_1655_io_out_0; // @[MUL.scala 104:13]
  assign m_1919_io_x3 = m_1652_io_out_1; // @[MUL.scala 105:13]
  assign m_1920_io_x1 = m_1656_io_s; // @[MUL.scala 252:21]
  assign m_1920_io_x2 = m_1653_io_cout; // @[MUL.scala 253:22]
  assign m_1920_io_x3 = m_1657_io_s; // @[MUL.scala 252:21]
  assign m_1921_io_x1 = m_1654_io_cout; // @[MUL.scala 253:22]
  assign m_1921_io_x2 = m_1658_io_out_0; // @[MUL.scala 104:13]
  assign m_1921_io_x3 = m_1655_io_out_1; // @[MUL.scala 105:13]
  assign m_1922_io_x1 = m_1659_io_s; // @[MUL.scala 252:21]
  assign m_1922_io_x2 = m_1656_io_cout; // @[MUL.scala 253:22]
  assign m_1922_io_x3 = m_1660_io_s; // @[MUL.scala 252:21]
  assign m_1923_io_x1 = m_1657_io_cout; // @[MUL.scala 253:22]
  assign m_1923_io_x2 = m_727_io_cout; // @[MUL.scala 253:22]
  assign m_1923_io_x3 = m_1658_io_out_1; // @[MUL.scala 105:13]
  assign m_1924_io_x1 = m_1661_io_s; // @[MUL.scala 252:21]
  assign m_1924_io_x2 = m_1659_io_cout; // @[MUL.scala 253:22]
  assign m_1924_io_x3 = m_1662_io_s; // @[MUL.scala 252:21]
  assign m_1925_io_in_0 = m_1660_io_cout; // @[MUL.scala 253:22]
  assign m_1925_io_in_1 = m_732_io_cout; // @[MUL.scala 253:22]
  assign m_1926_io_x1 = m_1663_io_s; // @[MUL.scala 252:21]
  assign m_1926_io_x2 = m_1661_io_cout; // @[MUL.scala 253:22]
  assign m_1926_io_x3 = m_1664_io_s; // @[MUL.scala 252:21]
  assign m_1927_io_in_0 = m_1662_io_cout; // @[MUL.scala 253:22]
  assign m_1927_io_in_1 = m_737_io_out_1; // @[MUL.scala 126:16]
  assign m_1928_io_x1 = m_1665_io_s; // @[MUL.scala 252:21]
  assign m_1928_io_x2 = m_1663_io_cout; // @[MUL.scala 253:22]
  assign m_1928_io_x3 = m_1666_io_s; // @[MUL.scala 252:21]
  assign m_1929_io_in_0 = m_1664_io_cout; // @[MUL.scala 253:22]
  assign m_1929_io_in_1 = m_742_io_out_1; // @[MUL.scala 126:16]
  assign m_1930_io_x1 = m_1667_io_s; // @[MUL.scala 252:21]
  assign m_1930_io_x2 = m_1665_io_cout; // @[MUL.scala 253:22]
  assign m_1930_io_x3 = m_1668_io_s; // @[MUL.scala 252:21]
  assign m_1931_io_x1 = m_1669_io_s; // @[MUL.scala 252:21]
  assign m_1931_io_x2 = m_1667_io_cout; // @[MUL.scala 253:22]
  assign m_1931_io_x3 = m_1670_io_s; // @[MUL.scala 252:21]
  assign m_1932_io_x1 = m_1671_io_s; // @[MUL.scala 252:21]
  assign m_1932_io_x2 = m_1669_io_cout; // @[MUL.scala 253:22]
  assign m_1932_io_x3 = m_1672_io_s; // @[MUL.scala 252:21]
  assign m_1933_io_x1 = m_1673_io_s; // @[MUL.scala 252:21]
  assign m_1933_io_x2 = m_1671_io_cout; // @[MUL.scala 253:22]
  assign m_1933_io_x3 = m_1674_io_s; // @[MUL.scala 252:21]
  assign m_1934_io_x1 = m_1675_io_s; // @[MUL.scala 252:21]
  assign m_1934_io_x2 = m_1673_io_cout; // @[MUL.scala 253:22]
  assign m_1934_io_x3 = m_1676_io_s; // @[MUL.scala 252:21]
  assign m_1935_io_x1 = m_1677_io_s; // @[MUL.scala 252:21]
  assign m_1935_io_x2 = m_1675_io_cout; // @[MUL.scala 253:22]
  assign m_1935_io_x3 = m_1678_io_s; // @[MUL.scala 252:21]
  assign m_1936_io_x1 = m_1679_io_s; // @[MUL.scala 252:21]
  assign m_1936_io_x2 = m_1677_io_cout; // @[MUL.scala 253:22]
  assign m_1936_io_x3 = m_1680_io_s; // @[MUL.scala 252:21]
  assign m_1937_io_x1 = m_1681_io_s; // @[MUL.scala 252:21]
  assign m_1937_io_x2 = m_1679_io_cout; // @[MUL.scala 253:22]
  assign m_1937_io_x3 = m_1305_io_cout; // @[MUL.scala 253:22]
  assign m_1938_io_x1 = m_1682_io_s; // @[MUL.scala 252:21]
  assign m_1938_io_x2 = m_1681_io_cout; // @[MUL.scala 253:22]
  assign m_1938_io_x3 = m_1307_io_cout; // @[MUL.scala 253:22]
  assign m_1939_io_x1 = m_1683_io_s; // @[MUL.scala 252:21]
  assign m_1939_io_x2 = m_1682_io_cout; // @[MUL.scala 253:22]
  assign m_1939_io_x3 = m_1309_io_cout; // @[MUL.scala 253:22]
  assign m_1940_io_x1 = m_1684_io_s; // @[MUL.scala 252:21]
  assign m_1940_io_x2 = m_1683_io_cout; // @[MUL.scala 253:22]
  assign m_1940_io_x3 = m_1311_io_cout; // @[MUL.scala 253:22]
  assign m_1941_io_x1 = m_1685_io_s; // @[MUL.scala 252:21]
  assign m_1941_io_x2 = m_1684_io_cout; // @[MUL.scala 253:22]
  assign m_1941_io_x3 = m_1313_io_cout; // @[MUL.scala 253:22]
  assign m_1942_io_x1 = m_1686_io_s; // @[MUL.scala 252:21]
  assign m_1942_io_x2 = m_1685_io_cout; // @[MUL.scala 253:22]
  assign m_1942_io_x3 = m_1315_io_cout; // @[MUL.scala 253:22]
  assign m_1943_io_x1 = m_1687_io_s; // @[MUL.scala 252:21]
  assign m_1943_io_x2 = m_1686_io_cout; // @[MUL.scala 253:22]
  assign m_1943_io_x3 = m_1317_io_out_1; // @[MUL.scala 105:13]
  assign m_1944_io_in_0 = m_1688_io_s; // @[MUL.scala 252:21]
  assign m_1944_io_in_1 = m_1687_io_cout; // @[MUL.scala 253:22]
  assign m_1945_io_in_0 = m_1689_io_s; // @[MUL.scala 252:21]
  assign m_1945_io_in_1 = m_1688_io_cout; // @[MUL.scala 253:22]
  assign m_1946_io_in_0 = m_1690_io_s; // @[MUL.scala 252:21]
  assign m_1946_io_in_1 = m_1689_io_cout; // @[MUL.scala 253:22]
  assign m_1947_io_in_0 = m_1691_io_s; // @[MUL.scala 252:21]
  assign m_1947_io_in_1 = m_1690_io_cout; // @[MUL.scala 253:22]
  assign m_1948_io_in_0 = m_1692_io_out_0; // @[MUL.scala 125:16]
  assign m_1948_io_in_1 = m_1691_io_cout; // @[MUL.scala 253:22]
  assign m_1949_io_in_0 = m_1693_io_out_0; // @[MUL.scala 125:16]
  assign m_1949_io_in_1 = m_1692_io_out_1; // @[MUL.scala 126:16]
  assign m_1950_io_in_0 = m_1694_io_out_0; // @[MUL.scala 125:16]
  assign m_1950_io_in_1 = m_1693_io_out_1; // @[MUL.scala 126:16]
  assign m_1951_io_in_0 = m_1695_io_out_0; // @[MUL.scala 125:16]
  assign m_1951_io_in_1 = m_1694_io_out_1; // @[MUL.scala 126:16]
  assign m_1952_io_in_0 = m_1696_io_out_0; // @[MUL.scala 125:16]
  assign m_1952_io_in_1 = m_1695_io_out_1; // @[MUL.scala 126:16]
  assign m_1953_io_in_0 = m_1697_io_out_0; // @[MUL.scala 125:16]
  assign m_1953_io_in_1 = m_1696_io_out_1; // @[MUL.scala 126:16]
  assign m_1954_io_in_0 = r_2312; // @[MUL.scala 125:16]
  assign m_1954_io_in_1 = r_2313; // @[MUL.scala 126:16]
  assign m_1955_io_in_0 = r_2314; // @[MUL.scala 125:16]
  assign m_1955_io_in_1 = r_2315; // @[MUL.scala 126:16]
  assign m_1956_io_in_0 = r_2316; // @[MUL.scala 125:16]
  assign m_1956_io_in_1 = r_2317; // @[MUL.scala 126:16]
  assign m_1957_io_in_0 = r_2318; // @[MUL.scala 125:16]
  assign m_1957_io_in_1 = r_2319; // @[MUL.scala 126:16]
  assign m_1958_io_in_0 = r_2320; // @[MUL.scala 125:16]
  assign m_1958_io_in_1 = r_2321; // @[MUL.scala 126:16]
  assign m_1959_io_in_0 = r_2322; // @[MUL.scala 125:16]
  assign m_1959_io_in_1 = r_2323; // @[MUL.scala 126:16]
  assign m_1960_io_in_0 = r_2324; // @[MUL.scala 125:16]
  assign m_1960_io_in_1 = r_2325; // @[MUL.scala 126:16]
  assign m_1961_io_in_0 = r_2326; // @[MUL.scala 125:16]
  assign m_1961_io_in_1 = r_2327; // @[MUL.scala 126:16]
  assign m_1962_io_in_0 = r_2328; // @[MUL.scala 125:16]
  assign m_1962_io_in_1 = r_2329; // @[MUL.scala 126:16]
  assign m_1963_io_in_0 = r_2330; // @[MUL.scala 125:16]
  assign m_1963_io_in_1 = r_2331; // @[MUL.scala 126:16]
  assign m_1964_io_in_0 = r_2332; // @[MUL.scala 125:16]
  assign m_1964_io_in_1 = r_2333; // @[MUL.scala 126:16]
  assign m_1965_io_in_0 = r_2334; // @[MUL.scala 125:16]
  assign m_1965_io_in_1 = r_2335; // @[MUL.scala 126:16]
  assign m_1966_io_in_0 = r_2336; // @[MUL.scala 125:16]
  assign m_1966_io_in_1 = r_2337; // @[MUL.scala 126:16]
  assign m_1967_io_x1 = r_2338; // @[MUL.scala 103:13]
  assign m_1967_io_x2 = r_2339; // @[MUL.scala 104:13]
  assign m_1967_io_x3 = r_2340; // @[MUL.scala 105:13]
  assign m_1968_io_x1 = r_2341; // @[MUL.scala 103:13]
  assign m_1968_io_x2 = r_2342; // @[MUL.scala 104:13]
  assign m_1968_io_x3 = r_2343; // @[MUL.scala 105:13]
  assign m_1969_io_x1 = r_2344; // @[MUL.scala 103:13]
  assign m_1969_io_x2 = r_2345; // @[MUL.scala 104:13]
  assign m_1969_io_x3 = r_2346; // @[MUL.scala 105:13]
  assign m_1970_io_x1 = r_2347; // @[MUL.scala 103:13]
  assign m_1970_io_x2 = r_2348; // @[MUL.scala 104:13]
  assign m_1970_io_x3 = r_2349; // @[MUL.scala 105:13]
  assign m_1971_io_x1 = r_2350; // @[MUL.scala 103:13]
  assign m_1971_io_x2 = r_2351; // @[MUL.scala 104:13]
  assign m_1971_io_x3 = r_2352; // @[MUL.scala 105:13]
  assign m_1972_io_x1 = r_2353; // @[MUL.scala 103:13]
  assign m_1972_io_x2 = r_2354; // @[MUL.scala 104:13]
  assign m_1972_io_x3 = r_2355; // @[MUL.scala 105:13]
  assign m_1973_io_x1 = r_2356; // @[MUL.scala 103:13]
  assign m_1973_io_x2 = r_2357; // @[MUL.scala 104:13]
  assign m_1973_io_x3 = r_2358; // @[MUL.scala 105:13]
  assign m_1974_io_x1 = r_2359; // @[MUL.scala 103:13]
  assign m_1974_io_x2 = r_2360; // @[MUL.scala 104:13]
  assign m_1974_io_x3 = r_2361; // @[MUL.scala 105:13]
  assign m_1975_io_x1 = r_2362; // @[MUL.scala 103:13]
  assign m_1975_io_x2 = r_2363; // @[MUL.scala 104:13]
  assign m_1975_io_x3 = r_2364; // @[MUL.scala 105:13]
  assign m_1976_io_x1 = r_2365; // @[MUL.scala 103:13]
  assign m_1976_io_x2 = r_2366; // @[MUL.scala 104:13]
  assign m_1976_io_x3 = r_2367; // @[MUL.scala 105:13]
  assign m_1977_io_x1 = r_2369; // @[MUL.scala 103:13]
  assign m_1977_io_x2 = r_2370; // @[MUL.scala 104:13]
  assign m_1977_io_x3 = r_2371; // @[MUL.scala 105:13]
  assign m_1978_io_x1 = r_2373; // @[MUL.scala 103:13]
  assign m_1978_io_x2 = r_2374; // @[MUL.scala 104:13]
  assign m_1978_io_x3 = r_2375; // @[MUL.scala 105:13]
  assign m_1979_io_x1 = r_2377; // @[MUL.scala 103:13]
  assign m_1979_io_x2 = r_2378; // @[MUL.scala 104:13]
  assign m_1979_io_x3 = r_2379; // @[MUL.scala 105:13]
  assign m_1980_io_x1 = r_2381; // @[MUL.scala 103:13]
  assign m_1980_io_x2 = r_2382; // @[MUL.scala 104:13]
  assign m_1980_io_x3 = r_2383; // @[MUL.scala 105:13]
  assign m_1981_io_x1 = r_2385; // @[MUL.scala 103:13]
  assign m_1981_io_x2 = r_2386; // @[MUL.scala 104:13]
  assign m_1981_io_x3 = r_2387; // @[MUL.scala 105:13]
  assign m_1982_io_x1 = r_2389; // @[MUL.scala 103:13]
  assign m_1982_io_x2 = r_2390; // @[MUL.scala 104:13]
  assign m_1982_io_x3 = r_2391; // @[MUL.scala 105:13]
  assign m_1983_io_x1 = r_2393; // @[MUL.scala 103:13]
  assign m_1983_io_x2 = r_2394; // @[MUL.scala 104:13]
  assign m_1983_io_x3 = r_2395; // @[MUL.scala 105:13]
  assign m_1984_io_x1 = r_2397; // @[MUL.scala 103:13]
  assign m_1984_io_x2 = r_2398; // @[MUL.scala 104:13]
  assign m_1984_io_x3 = r_2399; // @[MUL.scala 105:13]
  assign m_1985_io_x1 = r_2401; // @[MUL.scala 103:13]
  assign m_1985_io_x2 = r_2402; // @[MUL.scala 104:13]
  assign m_1985_io_x3 = r_2403; // @[MUL.scala 105:13]
  assign m_1986_io_x1 = r_2405; // @[MUL.scala 103:13]
  assign m_1986_io_x2 = r_2406; // @[MUL.scala 104:13]
  assign m_1986_io_x3 = r_2407; // @[MUL.scala 105:13]
  assign m_1987_io_x1 = r_2409; // @[MUL.scala 103:13]
  assign m_1987_io_x2 = r_2410; // @[MUL.scala 104:13]
  assign m_1987_io_x3 = r_2411; // @[MUL.scala 105:13]
  assign m_1988_io_x1 = r_2413; // @[MUL.scala 103:13]
  assign m_1988_io_x2 = r_2414; // @[MUL.scala 104:13]
  assign m_1988_io_x3 = r_2415; // @[MUL.scala 105:13]
  assign m_1989_io_in_0 = r_2416; // @[MUL.scala 125:16]
  assign m_1989_io_in_1 = r_2417; // @[MUL.scala 126:16]
  assign m_1990_io_x1 = r_2418; // @[MUL.scala 103:13]
  assign m_1990_io_x2 = r_2419; // @[MUL.scala 104:13]
  assign m_1990_io_x3 = r_2420; // @[MUL.scala 105:13]
  assign m_1991_io_in_0 = r_2421; // @[MUL.scala 125:16]
  assign m_1991_io_in_1 = r_2422; // @[MUL.scala 126:16]
  assign m_1992_io_x1 = r_2423; // @[MUL.scala 103:13]
  assign m_1992_io_x2 = r_2424; // @[MUL.scala 104:13]
  assign m_1992_io_x3 = r_2425; // @[MUL.scala 105:13]
  assign m_1993_io_in_0 = r_2426; // @[MUL.scala 125:16]
  assign m_1993_io_in_1 = r_2427; // @[MUL.scala 126:16]
  assign m_1994_io_x1 = r_2428; // @[MUL.scala 103:13]
  assign m_1994_io_x2 = r_2429; // @[MUL.scala 104:13]
  assign m_1994_io_x3 = r_2430; // @[MUL.scala 105:13]
  assign m_1995_io_in_0 = r_2431; // @[MUL.scala 125:16]
  assign m_1995_io_in_1 = r_2432; // @[MUL.scala 126:16]
  assign m_1996_io_x1 = r_2433; // @[MUL.scala 103:13]
  assign m_1996_io_x2 = r_2434; // @[MUL.scala 104:13]
  assign m_1996_io_x3 = r_2435; // @[MUL.scala 105:13]
  assign m_1997_io_in_0 = r_2436; // @[MUL.scala 125:16]
  assign m_1997_io_in_1 = r_2437; // @[MUL.scala 126:16]
  assign m_1998_io_x1 = r_2438; // @[MUL.scala 103:13]
  assign m_1998_io_x2 = r_2439; // @[MUL.scala 104:13]
  assign m_1998_io_x3 = r_2440; // @[MUL.scala 105:13]
  assign m_1999_io_in_0 = r_2441; // @[MUL.scala 125:16]
  assign m_1999_io_in_1 = r_2442; // @[MUL.scala 126:16]
  assign m_2000_io_x1 = r_2443; // @[MUL.scala 103:13]
  assign m_2000_io_x2 = r_2444; // @[MUL.scala 104:13]
  assign m_2000_io_x3 = r_2445; // @[MUL.scala 105:13]
  assign m_2001_io_in_0 = r_2446; // @[MUL.scala 125:16]
  assign m_2001_io_in_1 = r_2447; // @[MUL.scala 126:16]
  assign m_2002_io_x1 = r_2448; // @[MUL.scala 103:13]
  assign m_2002_io_x2 = r_2449; // @[MUL.scala 104:13]
  assign m_2002_io_x3 = r_2450; // @[MUL.scala 105:13]
  assign m_2003_io_x1 = r_2451; // @[MUL.scala 103:13]
  assign m_2003_io_x2 = r_2452; // @[MUL.scala 104:13]
  assign m_2003_io_x3 = r_2453; // @[MUL.scala 105:13]
  assign m_2004_io_x1 = r_2454; // @[MUL.scala 103:13]
  assign m_2004_io_x2 = r_2455; // @[MUL.scala 104:13]
  assign m_2004_io_x3 = r_2456; // @[MUL.scala 105:13]
  assign m_2005_io_x1 = r_2457; // @[MUL.scala 103:13]
  assign m_2005_io_x2 = r_2458; // @[MUL.scala 104:13]
  assign m_2005_io_x3 = r_2459; // @[MUL.scala 105:13]
  assign m_2006_io_x1 = r_2460; // @[MUL.scala 103:13]
  assign m_2006_io_x2 = r_2461; // @[MUL.scala 104:13]
  assign m_2006_io_x3 = r_2462; // @[MUL.scala 105:13]
  assign m_2007_io_x1 = r_2463; // @[MUL.scala 103:13]
  assign m_2007_io_x2 = r_2464; // @[MUL.scala 104:13]
  assign m_2007_io_x3 = r_2465; // @[MUL.scala 105:13]
  assign m_2008_io_x1 = r_2466; // @[MUL.scala 103:13]
  assign m_2008_io_x2 = r_2467; // @[MUL.scala 104:13]
  assign m_2008_io_x3 = r_2468; // @[MUL.scala 105:13]
  assign m_2009_io_x1 = r_2469; // @[MUL.scala 103:13]
  assign m_2009_io_x2 = r_2470; // @[MUL.scala 104:13]
  assign m_2009_io_x3 = r_2471; // @[MUL.scala 105:13]
  assign m_2010_io_x1 = r_2472; // @[MUL.scala 103:13]
  assign m_2010_io_x2 = r_2473; // @[MUL.scala 104:13]
  assign m_2010_io_x3 = r_2474; // @[MUL.scala 105:13]
  assign m_2011_io_x1 = r_2475; // @[MUL.scala 103:13]
  assign m_2011_io_x2 = r_2476; // @[MUL.scala 104:13]
  assign m_2011_io_x3 = r_2477; // @[MUL.scala 105:13]
  assign m_2012_io_x1 = r_2478; // @[MUL.scala 103:13]
  assign m_2012_io_x2 = r_2479; // @[MUL.scala 104:13]
  assign m_2012_io_x3 = r_2480; // @[MUL.scala 105:13]
  assign m_2013_io_x1 = r_2481; // @[MUL.scala 103:13]
  assign m_2013_io_x2 = r_2482; // @[MUL.scala 104:13]
  assign m_2013_io_x3 = r_2483; // @[MUL.scala 105:13]
  assign m_2014_io_x1 = r_2484; // @[MUL.scala 103:13]
  assign m_2014_io_x2 = r_2485; // @[MUL.scala 104:13]
  assign m_2014_io_x3 = r_2486; // @[MUL.scala 105:13]
  assign m_2015_io_x1 = r_2487; // @[MUL.scala 103:13]
  assign m_2015_io_x2 = r_2488; // @[MUL.scala 104:13]
  assign m_2015_io_x3 = r_2489; // @[MUL.scala 105:13]
  assign m_2016_io_x1 = r_2490; // @[MUL.scala 103:13]
  assign m_2016_io_x2 = r_2491; // @[MUL.scala 104:13]
  assign m_2016_io_x3 = r_2492; // @[MUL.scala 105:13]
  assign m_2017_io_x1 = r_2493; // @[MUL.scala 103:13]
  assign m_2017_io_x2 = r_2494; // @[MUL.scala 104:13]
  assign m_2017_io_x3 = r_2495; // @[MUL.scala 105:13]
  assign m_2018_io_x1 = r_2496; // @[MUL.scala 103:13]
  assign m_2018_io_x2 = r_2497; // @[MUL.scala 104:13]
  assign m_2018_io_x3 = r_2498; // @[MUL.scala 105:13]
  assign m_2019_io_x1 = r_2499; // @[MUL.scala 103:13]
  assign m_2019_io_x2 = r_2500; // @[MUL.scala 104:13]
  assign m_2019_io_x3 = r_2501; // @[MUL.scala 105:13]
  assign m_2020_io_x1 = r_2502; // @[MUL.scala 103:13]
  assign m_2020_io_x2 = r_2503; // @[MUL.scala 104:13]
  assign m_2020_io_x3 = r_2504; // @[MUL.scala 105:13]
  assign m_2021_io_x1 = r_2505; // @[MUL.scala 103:13]
  assign m_2021_io_x2 = r_2506; // @[MUL.scala 104:13]
  assign m_2021_io_x3 = r_2507; // @[MUL.scala 105:13]
  assign m_2022_io_x1 = r_2508; // @[MUL.scala 103:13]
  assign m_2022_io_x2 = r_2509; // @[MUL.scala 104:13]
  assign m_2022_io_x3 = r_2510; // @[MUL.scala 105:13]
  assign m_2023_io_x1 = r_2511; // @[MUL.scala 103:13]
  assign m_2023_io_x2 = r_2512; // @[MUL.scala 104:13]
  assign m_2023_io_x3 = r_2513; // @[MUL.scala 105:13]
  assign m_2024_io_x1 = r_2514; // @[MUL.scala 103:13]
  assign m_2024_io_x2 = r_2515; // @[MUL.scala 104:13]
  assign m_2024_io_x3 = r_2516; // @[MUL.scala 105:13]
  assign m_2025_io_x1 = r_2517; // @[MUL.scala 103:13]
  assign m_2025_io_x2 = r_2518; // @[MUL.scala 104:13]
  assign m_2025_io_x3 = r_2519; // @[MUL.scala 105:13]
  assign m_2026_io_x1 = r_2520; // @[MUL.scala 103:13]
  assign m_2026_io_x2 = r_2521; // @[MUL.scala 104:13]
  assign m_2026_io_x3 = r_2522; // @[MUL.scala 105:13]
  assign m_2027_io_x1 = r_2523; // @[MUL.scala 103:13]
  assign m_2027_io_x2 = r_2524; // @[MUL.scala 104:13]
  assign m_2027_io_x3 = r_2525; // @[MUL.scala 105:13]
  assign m_2028_io_x1 = r_2527; // @[MUL.scala 103:13]
  assign m_2028_io_x2 = r_2528; // @[MUL.scala 104:13]
  assign m_2028_io_x3 = r_2529; // @[MUL.scala 105:13]
  assign m_2029_io_x1 = r_2530; // @[MUL.scala 103:13]
  assign m_2029_io_x2 = r_2531; // @[MUL.scala 104:13]
  assign m_2029_io_x3 = r_2532; // @[MUL.scala 105:13]
  assign m_2030_io_x1 = r_2534; // @[MUL.scala 103:13]
  assign m_2030_io_x2 = r_2535; // @[MUL.scala 104:13]
  assign m_2030_io_x3 = r_2536; // @[MUL.scala 105:13]
  assign m_2031_io_x1 = r_2537; // @[MUL.scala 103:13]
  assign m_2031_io_x2 = r_2538; // @[MUL.scala 104:13]
  assign m_2031_io_x3 = r_2539; // @[MUL.scala 105:13]
  assign m_2032_io_x1 = r_2541; // @[MUL.scala 103:13]
  assign m_2032_io_x2 = r_2542; // @[MUL.scala 104:13]
  assign m_2032_io_x3 = r_2543; // @[MUL.scala 105:13]
  assign m_2033_io_x1 = r_2544; // @[MUL.scala 103:13]
  assign m_2033_io_x2 = r_2545; // @[MUL.scala 104:13]
  assign m_2033_io_x3 = r_2546; // @[MUL.scala 105:13]
  assign m_2034_io_x1 = r_2548; // @[MUL.scala 103:13]
  assign m_2034_io_x2 = r_2549; // @[MUL.scala 104:13]
  assign m_2034_io_x3 = r_2550; // @[MUL.scala 105:13]
  assign m_2035_io_x1 = r_2551; // @[MUL.scala 103:13]
  assign m_2035_io_x2 = r_2552; // @[MUL.scala 104:13]
  assign m_2035_io_x3 = r_2553; // @[MUL.scala 105:13]
  assign m_2036_io_x1 = r_2555; // @[MUL.scala 103:13]
  assign m_2036_io_x2 = r_2556; // @[MUL.scala 104:13]
  assign m_2036_io_x3 = r_2557; // @[MUL.scala 105:13]
  assign m_2037_io_x1 = r_2558; // @[MUL.scala 103:13]
  assign m_2037_io_x2 = r_2559; // @[MUL.scala 104:13]
  assign m_2037_io_x3 = r_2560; // @[MUL.scala 105:13]
  assign m_2038_io_x1 = r_2562; // @[MUL.scala 103:13]
  assign m_2038_io_x2 = r_2563; // @[MUL.scala 104:13]
  assign m_2038_io_x3 = r_2564; // @[MUL.scala 105:13]
  assign m_2039_io_x1 = r_2565; // @[MUL.scala 103:13]
  assign m_2039_io_x2 = r_2566; // @[MUL.scala 104:13]
  assign m_2039_io_x3 = r_2567; // @[MUL.scala 105:13]
  assign m_2040_io_x1 = r_2569; // @[MUL.scala 103:13]
  assign m_2040_io_x2 = r_2570; // @[MUL.scala 104:13]
  assign m_2040_io_x3 = r_2571; // @[MUL.scala 105:13]
  assign m_2041_io_x1 = r_2572; // @[MUL.scala 103:13]
  assign m_2041_io_x2 = r_2573; // @[MUL.scala 104:13]
  assign m_2041_io_x3 = r_2574; // @[MUL.scala 105:13]
  assign m_2042_io_x1 = r_2576; // @[MUL.scala 103:13]
  assign m_2042_io_x2 = r_2577; // @[MUL.scala 104:13]
  assign m_2042_io_x3 = r_2578; // @[MUL.scala 105:13]
  assign m_2043_io_x1 = r_2579; // @[MUL.scala 103:13]
  assign m_2043_io_x2 = r_2580; // @[MUL.scala 104:13]
  assign m_2043_io_x3 = r_2581; // @[MUL.scala 105:13]
  assign m_2044_io_x1 = r_2583; // @[MUL.scala 103:13]
  assign m_2044_io_x2 = r_2584; // @[MUL.scala 104:13]
  assign m_2044_io_x3 = r_2585; // @[MUL.scala 105:13]
  assign m_2045_io_x1 = r_2586; // @[MUL.scala 103:13]
  assign m_2045_io_x2 = r_2587; // @[MUL.scala 104:13]
  assign m_2045_io_x3 = r_2588; // @[MUL.scala 105:13]
  assign m_2046_io_x1 = r_2590; // @[MUL.scala 103:13]
  assign m_2046_io_x2 = r_2591; // @[MUL.scala 104:13]
  assign m_2046_io_x3 = r_2592; // @[MUL.scala 105:13]
  assign m_2047_io_x1 = r_2593; // @[MUL.scala 103:13]
  assign m_2047_io_x2 = r_2594; // @[MUL.scala 104:13]
  assign m_2047_io_x3 = r_2595; // @[MUL.scala 105:13]
  assign m_2048_io_x1 = r_2597; // @[MUL.scala 103:13]
  assign m_2048_io_x2 = r_2598; // @[MUL.scala 104:13]
  assign m_2048_io_x3 = r_2599; // @[MUL.scala 105:13]
  assign m_2049_io_x1 = r_2600; // @[MUL.scala 103:13]
  assign m_2049_io_x2 = r_2601; // @[MUL.scala 104:13]
  assign m_2049_io_x3 = r_2602; // @[MUL.scala 105:13]
  assign m_2050_io_x1 = r_2604; // @[MUL.scala 103:13]
  assign m_2050_io_x2 = r_2605; // @[MUL.scala 104:13]
  assign m_2050_io_x3 = r_2606; // @[MUL.scala 105:13]
  assign m_2051_io_x1 = r_2607; // @[MUL.scala 103:13]
  assign m_2051_io_x2 = r_2608; // @[MUL.scala 104:13]
  assign m_2051_io_x3 = r_2609; // @[MUL.scala 105:13]
  assign m_2052_io_x1 = r_2611; // @[MUL.scala 103:13]
  assign m_2052_io_x2 = r_2612; // @[MUL.scala 104:13]
  assign m_2052_io_x3 = r_2613; // @[MUL.scala 105:13]
  assign m_2053_io_x1 = r_2614; // @[MUL.scala 103:13]
  assign m_2053_io_x2 = r_2615; // @[MUL.scala 104:13]
  assign m_2053_io_x3 = r_2616; // @[MUL.scala 105:13]
  assign m_2054_io_x1 = r_2618; // @[MUL.scala 103:13]
  assign m_2054_io_x2 = r_2619; // @[MUL.scala 104:13]
  assign m_2054_io_x3 = r_2620; // @[MUL.scala 105:13]
  assign m_2055_io_x1 = r_2621; // @[MUL.scala 103:13]
  assign m_2055_io_x2 = r_2622; // @[MUL.scala 104:13]
  assign m_2055_io_x3 = r_2623; // @[MUL.scala 105:13]
  assign m_2056_io_x1 = r_2625; // @[MUL.scala 103:13]
  assign m_2056_io_x2 = r_2626; // @[MUL.scala 104:13]
  assign m_2056_io_x3 = r_2627; // @[MUL.scala 105:13]
  assign m_2057_io_x1 = r_2628; // @[MUL.scala 103:13]
  assign m_2057_io_x2 = r_2629; // @[MUL.scala 104:13]
  assign m_2057_io_x3 = r_2630; // @[MUL.scala 105:13]
  assign m_2058_io_x1 = r_2632; // @[MUL.scala 103:13]
  assign m_2058_io_x2 = r_2633; // @[MUL.scala 104:13]
  assign m_2058_io_x3 = r_2634; // @[MUL.scala 105:13]
  assign m_2059_io_x1 = r_2635; // @[MUL.scala 103:13]
  assign m_2059_io_x2 = r_2636; // @[MUL.scala 104:13]
  assign m_2059_io_x3 = r_2637; // @[MUL.scala 105:13]
  assign m_2060_io_x1 = r_2639; // @[MUL.scala 103:13]
  assign m_2060_io_x2 = r_2640; // @[MUL.scala 104:13]
  assign m_2060_io_x3 = r_2641; // @[MUL.scala 105:13]
  assign m_2061_io_x1 = r_2642; // @[MUL.scala 103:13]
  assign m_2061_io_x2 = r_2643; // @[MUL.scala 104:13]
  assign m_2061_io_x3 = r_2644; // @[MUL.scala 105:13]
  assign m_2062_io_x1 = r_2646; // @[MUL.scala 103:13]
  assign m_2062_io_x2 = r_2647; // @[MUL.scala 104:13]
  assign m_2062_io_x3 = r_2648; // @[MUL.scala 105:13]
  assign m_2063_io_x1 = r_2649; // @[MUL.scala 103:13]
  assign m_2063_io_x2 = r_2650; // @[MUL.scala 104:13]
  assign m_2063_io_x3 = r_2651; // @[MUL.scala 105:13]
  assign m_2064_io_x1 = r_2653; // @[MUL.scala 103:13]
  assign m_2064_io_x2 = r_2654; // @[MUL.scala 104:13]
  assign m_2064_io_x3 = r_2655; // @[MUL.scala 105:13]
  assign m_2065_io_x1 = r_2656; // @[MUL.scala 103:13]
  assign m_2065_io_x2 = r_2657; // @[MUL.scala 104:13]
  assign m_2065_io_x3 = r_2658; // @[MUL.scala 105:13]
  assign m_2066_io_x1 = r_2660; // @[MUL.scala 103:13]
  assign m_2066_io_x2 = r_2661; // @[MUL.scala 104:13]
  assign m_2066_io_x3 = r_2662; // @[MUL.scala 105:13]
  assign m_2067_io_x1 = r_2663; // @[MUL.scala 103:13]
  assign m_2067_io_x2 = r_2664; // @[MUL.scala 104:13]
  assign m_2067_io_x3 = r_2665; // @[MUL.scala 105:13]
  assign m_2068_io_x1 = r_2667; // @[MUL.scala 103:13]
  assign m_2068_io_x2 = r_2668; // @[MUL.scala 104:13]
  assign m_2068_io_x3 = r_2669; // @[MUL.scala 105:13]
  assign m_2069_io_x1 = r_2670; // @[MUL.scala 103:13]
  assign m_2069_io_x2 = r_2671; // @[MUL.scala 104:13]
  assign m_2069_io_x3 = r_2672; // @[MUL.scala 105:13]
  assign m_2070_io_x1 = r_2673; // @[MUL.scala 103:13]
  assign m_2070_io_x2 = r_2674; // @[MUL.scala 104:13]
  assign m_2070_io_x3 = r_2675; // @[MUL.scala 105:13]
  assign m_2071_io_x1 = r_2676; // @[MUL.scala 103:13]
  assign m_2071_io_x2 = r_2677; // @[MUL.scala 104:13]
  assign m_2071_io_x3 = r_2678; // @[MUL.scala 105:13]
  assign m_2072_io_x1 = r_2679; // @[MUL.scala 103:13]
  assign m_2072_io_x2 = r_2680; // @[MUL.scala 104:13]
  assign m_2072_io_x3 = r_2681; // @[MUL.scala 105:13]
  assign m_2073_io_x1 = r_2682; // @[MUL.scala 103:13]
  assign m_2073_io_x2 = r_2683; // @[MUL.scala 104:13]
  assign m_2073_io_x3 = r_2684; // @[MUL.scala 105:13]
  assign m_2074_io_x1 = r_2685; // @[MUL.scala 103:13]
  assign m_2074_io_x2 = r_2686; // @[MUL.scala 104:13]
  assign m_2074_io_x3 = r_2687; // @[MUL.scala 105:13]
  assign m_2075_io_x1 = r_2688; // @[MUL.scala 103:13]
  assign m_2075_io_x2 = r_2689; // @[MUL.scala 104:13]
  assign m_2075_io_x3 = r_2690; // @[MUL.scala 105:13]
  assign m_2076_io_x1 = r_2691; // @[MUL.scala 103:13]
  assign m_2076_io_x2 = r_2692; // @[MUL.scala 104:13]
  assign m_2076_io_x3 = r_2693; // @[MUL.scala 105:13]
  assign m_2077_io_x1 = r_2694; // @[MUL.scala 103:13]
  assign m_2077_io_x2 = r_2695; // @[MUL.scala 104:13]
  assign m_2077_io_x3 = r_2696; // @[MUL.scala 105:13]
  assign m_2078_io_x1 = r_2697; // @[MUL.scala 103:13]
  assign m_2078_io_x2 = r_2698; // @[MUL.scala 104:13]
  assign m_2078_io_x3 = r_2699; // @[MUL.scala 105:13]
  assign m_2079_io_x1 = r_2700; // @[MUL.scala 103:13]
  assign m_2079_io_x2 = r_2701; // @[MUL.scala 104:13]
  assign m_2079_io_x3 = r_2702; // @[MUL.scala 105:13]
  assign m_2080_io_x1 = r_2703; // @[MUL.scala 103:13]
  assign m_2080_io_x2 = r_2704; // @[MUL.scala 104:13]
  assign m_2080_io_x3 = r_2705; // @[MUL.scala 105:13]
  assign m_2081_io_x1 = r_2706; // @[MUL.scala 103:13]
  assign m_2081_io_x2 = r_2707; // @[MUL.scala 104:13]
  assign m_2081_io_x3 = r_2708; // @[MUL.scala 105:13]
  assign m_2082_io_x1 = r_2709; // @[MUL.scala 103:13]
  assign m_2082_io_x2 = r_2710; // @[MUL.scala 104:13]
  assign m_2082_io_x3 = r_2711; // @[MUL.scala 105:13]
  assign m_2083_io_x1 = r_2712; // @[MUL.scala 103:13]
  assign m_2083_io_x2 = r_2713; // @[MUL.scala 104:13]
  assign m_2083_io_x3 = r_2714; // @[MUL.scala 105:13]
  assign m_2084_io_x1 = r_2715; // @[MUL.scala 103:13]
  assign m_2084_io_x2 = r_2716; // @[MUL.scala 104:13]
  assign m_2084_io_x3 = r_2717; // @[MUL.scala 105:13]
  assign m_2085_io_x1 = r_2718; // @[MUL.scala 103:13]
  assign m_2085_io_x2 = r_2719; // @[MUL.scala 104:13]
  assign m_2085_io_x3 = r_2720; // @[MUL.scala 105:13]
  assign m_2086_io_x1 = r_2721; // @[MUL.scala 103:13]
  assign m_2086_io_x2 = r_2722; // @[MUL.scala 104:13]
  assign m_2086_io_x3 = r_2723; // @[MUL.scala 105:13]
  assign m_2087_io_x1 = r_2724; // @[MUL.scala 103:13]
  assign m_2087_io_x2 = r_2725; // @[MUL.scala 104:13]
  assign m_2087_io_x3 = r_2726; // @[MUL.scala 105:13]
  assign m_2088_io_x1 = r_2727; // @[MUL.scala 103:13]
  assign m_2088_io_x2 = r_2728; // @[MUL.scala 104:13]
  assign m_2088_io_x3 = r_2729; // @[MUL.scala 105:13]
  assign m_2089_io_x1 = r_2730; // @[MUL.scala 103:13]
  assign m_2089_io_x2 = r_2731; // @[MUL.scala 104:13]
  assign m_2089_io_x3 = r_2732; // @[MUL.scala 105:13]
  assign m_2090_io_x1 = r_2733; // @[MUL.scala 103:13]
  assign m_2090_io_x2 = r_2734; // @[MUL.scala 104:13]
  assign m_2090_io_x3 = r_2735; // @[MUL.scala 105:13]
  assign m_2091_io_x1 = r_2736; // @[MUL.scala 103:13]
  assign m_2091_io_x2 = r_2737; // @[MUL.scala 104:13]
  assign m_2091_io_x3 = r_2738; // @[MUL.scala 105:13]
  assign m_2092_io_x1 = r_2739; // @[MUL.scala 103:13]
  assign m_2092_io_x2 = r_2740; // @[MUL.scala 104:13]
  assign m_2092_io_x3 = r_2741; // @[MUL.scala 105:13]
  assign m_2093_io_x1 = r_2742; // @[MUL.scala 103:13]
  assign m_2093_io_x2 = r_2743; // @[MUL.scala 104:13]
  assign m_2093_io_x3 = r_2744; // @[MUL.scala 105:13]
  assign m_2094_io_x1 = r_2745; // @[MUL.scala 103:13]
  assign m_2094_io_x2 = r_2746; // @[MUL.scala 104:13]
  assign m_2094_io_x3 = r_2747; // @[MUL.scala 105:13]
  assign m_2095_io_in_0 = r_2748; // @[MUL.scala 125:16]
  assign m_2095_io_in_1 = r_2749; // @[MUL.scala 126:16]
  assign m_2096_io_x1 = r_2750; // @[MUL.scala 103:13]
  assign m_2096_io_x2 = r_2751; // @[MUL.scala 104:13]
  assign m_2096_io_x3 = r_2752; // @[MUL.scala 105:13]
  assign m_2097_io_in_0 = r_2753; // @[MUL.scala 125:16]
  assign m_2097_io_in_1 = r_2754; // @[MUL.scala 126:16]
  assign m_2098_io_x1 = r_2755; // @[MUL.scala 103:13]
  assign m_2098_io_x2 = r_2756; // @[MUL.scala 104:13]
  assign m_2098_io_x3 = r_2757; // @[MUL.scala 105:13]
  assign m_2099_io_in_0 = r_2758; // @[MUL.scala 125:16]
  assign m_2099_io_in_1 = r_2759; // @[MUL.scala 126:16]
  assign m_2100_io_x1 = r_2760; // @[MUL.scala 103:13]
  assign m_2100_io_x2 = r_2761; // @[MUL.scala 104:13]
  assign m_2100_io_x3 = r_2762; // @[MUL.scala 105:13]
  assign m_2101_io_in_0 = r_2763; // @[MUL.scala 125:16]
  assign m_2101_io_in_1 = r_2764; // @[MUL.scala 126:16]
  assign m_2102_io_x1 = r_2765; // @[MUL.scala 103:13]
  assign m_2102_io_x2 = r_2766; // @[MUL.scala 104:13]
  assign m_2102_io_x3 = r_2767; // @[MUL.scala 105:13]
  assign m_2103_io_in_0 = r_2768; // @[MUL.scala 125:16]
  assign m_2103_io_in_1 = r_2769; // @[MUL.scala 126:16]
  assign m_2104_io_x1 = r_2770; // @[MUL.scala 103:13]
  assign m_2104_io_x2 = r_2771; // @[MUL.scala 104:13]
  assign m_2104_io_x3 = r_2772; // @[MUL.scala 105:13]
  assign m_2105_io_x1 = r_2774; // @[MUL.scala 103:13]
  assign m_2105_io_x2 = r_2775; // @[MUL.scala 104:13]
  assign m_2105_io_x3 = r_2776; // @[MUL.scala 105:13]
  assign m_2106_io_x1 = r_2778; // @[MUL.scala 103:13]
  assign m_2106_io_x2 = r_2779; // @[MUL.scala 104:13]
  assign m_2106_io_x3 = r_2780; // @[MUL.scala 105:13]
  assign m_2107_io_x1 = r_2782; // @[MUL.scala 103:13]
  assign m_2107_io_x2 = r_2783; // @[MUL.scala 104:13]
  assign m_2107_io_x3 = r_2784; // @[MUL.scala 105:13]
  assign m_2108_io_x1 = r_2786; // @[MUL.scala 103:13]
  assign m_2108_io_x2 = r_2787; // @[MUL.scala 104:13]
  assign m_2108_io_x3 = r_2788; // @[MUL.scala 105:13]
  assign m_2109_io_x1 = r_2790; // @[MUL.scala 103:13]
  assign m_2109_io_x2 = r_2791; // @[MUL.scala 104:13]
  assign m_2109_io_x3 = r_2792; // @[MUL.scala 105:13]
  assign m_2110_io_x1 = r_2794; // @[MUL.scala 103:13]
  assign m_2110_io_x2 = r_2795; // @[MUL.scala 104:13]
  assign m_2110_io_x3 = r_2796; // @[MUL.scala 105:13]
  assign m_2111_io_x1 = r_2798; // @[MUL.scala 103:13]
  assign m_2111_io_x2 = r_2799; // @[MUL.scala 104:13]
  assign m_2111_io_x3 = r_2800; // @[MUL.scala 105:13]
  assign m_2112_io_x1 = r_2802; // @[MUL.scala 103:13]
  assign m_2112_io_x2 = r_2803; // @[MUL.scala 104:13]
  assign m_2112_io_x3 = r_2804; // @[MUL.scala 105:13]
  assign m_2113_io_x1 = r_2806; // @[MUL.scala 103:13]
  assign m_2113_io_x2 = r_2807; // @[MUL.scala 104:13]
  assign m_2113_io_x3 = r_2808; // @[MUL.scala 105:13]
  assign m_2114_io_x1 = r_2810; // @[MUL.scala 103:13]
  assign m_2114_io_x2 = r_2811; // @[MUL.scala 104:13]
  assign m_2114_io_x3 = r_2812; // @[MUL.scala 105:13]
  assign m_2115_io_x1 = r_2814; // @[MUL.scala 103:13]
  assign m_2115_io_x2 = r_2815; // @[MUL.scala 104:13]
  assign m_2115_io_x3 = r_2816; // @[MUL.scala 105:13]
  assign m_2116_io_x1 = r_2818; // @[MUL.scala 103:13]
  assign m_2116_io_x2 = r_2819; // @[MUL.scala 104:13]
  assign m_2116_io_x3 = r_2820; // @[MUL.scala 105:13]
  assign m_2117_io_x1 = r_2821; // @[MUL.scala 103:13]
  assign m_2117_io_x2 = r_2822; // @[MUL.scala 104:13]
  assign m_2117_io_x3 = r_2823; // @[MUL.scala 105:13]
  assign m_2118_io_x1 = r_2824; // @[MUL.scala 103:13]
  assign m_2118_io_x2 = r_2825; // @[MUL.scala 104:13]
  assign m_2118_io_x3 = r_2826; // @[MUL.scala 105:13]
  assign m_2119_io_x1 = r_2827; // @[MUL.scala 103:13]
  assign m_2119_io_x2 = r_2828; // @[MUL.scala 104:13]
  assign m_2119_io_x3 = r_2829; // @[MUL.scala 105:13]
  assign m_2120_io_x1 = r_2830; // @[MUL.scala 103:13]
  assign m_2120_io_x2 = r_2831; // @[MUL.scala 104:13]
  assign m_2120_io_x3 = r_2832; // @[MUL.scala 105:13]
  assign m_2121_io_x1 = r_2833; // @[MUL.scala 103:13]
  assign m_2121_io_x2 = r_2834; // @[MUL.scala 104:13]
  assign m_2121_io_x3 = r_2835; // @[MUL.scala 105:13]
  assign m_2122_io_x1 = r_2836; // @[MUL.scala 103:13]
  assign m_2122_io_x2 = r_2837; // @[MUL.scala 104:13]
  assign m_2122_io_x3 = r_2838; // @[MUL.scala 105:13]
  assign m_2123_io_in_0 = r_2839; // @[MUL.scala 125:16]
  assign m_2123_io_in_1 = r_2840; // @[MUL.scala 126:16]
  assign m_2124_io_in_0 = r_2841; // @[MUL.scala 125:16]
  assign m_2124_io_in_1 = r_2842; // @[MUL.scala 126:16]
  assign m_2125_io_in_0 = r_2843; // @[MUL.scala 125:16]
  assign m_2125_io_in_1 = r_2844; // @[MUL.scala 126:16]
  assign m_2126_io_in_0 = r_2845; // @[MUL.scala 125:16]
  assign m_2126_io_in_1 = r_2846; // @[MUL.scala 126:16]
  assign m_2127_io_in_0 = r_2847; // @[MUL.scala 125:16]
  assign m_2127_io_in_1 = r_2848; // @[MUL.scala 126:16]
  assign m_2128_io_in_0 = r_2849; // @[MUL.scala 125:16]
  assign m_2128_io_in_1 = r_2850; // @[MUL.scala 126:16]
  assign m_2129_io_in_0 = r_2851; // @[MUL.scala 125:16]
  assign m_2129_io_in_1 = r_2852; // @[MUL.scala 126:16]
  assign m_2130_io_in_0 = r_2853; // @[MUL.scala 125:16]
  assign m_2130_io_in_1 = r_2854; // @[MUL.scala 126:16]
  assign m_2131_io_in_0 = r_2855; // @[MUL.scala 125:16]
  assign m_2131_io_in_1 = r_2856; // @[MUL.scala 126:16]
  assign m_2132_io_in_0 = r_2857; // @[MUL.scala 125:16]
  assign m_2132_io_in_1 = r_2858; // @[MUL.scala 126:16]
  assign m_2133_io_in_0 = r_2859; // @[MUL.scala 125:16]
  assign m_2133_io_in_1 = r_2860; // @[MUL.scala 126:16]
  assign m_2134_io_in_0 = r_2861; // @[MUL.scala 125:16]
  assign m_2134_io_in_1 = r_2862; // @[MUL.scala 126:16]
  assign m_2135_io_in_0 = r_2863; // @[MUL.scala 125:16]
  assign m_2135_io_in_1 = r_2864; // @[MUL.scala 126:16]
  assign m_2136_io_in_0 = r_2865; // @[MUL.scala 125:16]
  assign m_2136_io_in_1 = r_2866; // @[MUL.scala 126:16]
  assign m_2137_io_in_0 = r_2867; // @[MUL.scala 125:16]
  assign m_2137_io_in_1 = r_2868; // @[MUL.scala 126:16]
  assign m_2138_io_in_0 = r_2869; // @[MUL.scala 125:16]
  assign m_2138_io_in_1 = r_2870; // @[MUL.scala 126:16]
  assign m_2139_io_in_0 = m_1955_io_out_0; // @[MUL.scala 125:16]
  assign m_2139_io_in_1 = m_1954_io_out_1; // @[MUL.scala 126:16]
  assign m_2140_io_in_0 = m_1956_io_out_0; // @[MUL.scala 125:16]
  assign m_2140_io_in_1 = m_1955_io_out_1; // @[MUL.scala 126:16]
  assign m_2141_io_in_0 = m_1957_io_out_0; // @[MUL.scala 125:16]
  assign m_2141_io_in_1 = m_1956_io_out_1; // @[MUL.scala 126:16]
  assign m_2142_io_in_0 = m_1958_io_out_0; // @[MUL.scala 125:16]
  assign m_2142_io_in_1 = m_1957_io_out_1; // @[MUL.scala 126:16]
  assign m_2143_io_in_0 = m_1959_io_out_0; // @[MUL.scala 125:16]
  assign m_2143_io_in_1 = m_1958_io_out_1; // @[MUL.scala 126:16]
  assign m_2144_io_in_0 = m_1960_io_out_0; // @[MUL.scala 125:16]
  assign m_2144_io_in_1 = m_1959_io_out_1; // @[MUL.scala 126:16]
  assign m_2145_io_in_0 = m_1961_io_out_0; // @[MUL.scala 125:16]
  assign m_2145_io_in_1 = m_1960_io_out_1; // @[MUL.scala 126:16]
  assign m_2146_io_in_0 = m_1962_io_out_0; // @[MUL.scala 125:16]
  assign m_2146_io_in_1 = m_1961_io_out_1; // @[MUL.scala 126:16]
  assign m_2147_io_in_0 = m_1963_io_out_0; // @[MUL.scala 125:16]
  assign m_2147_io_in_1 = m_1962_io_out_1; // @[MUL.scala 126:16]
  assign m_2148_io_in_0 = m_1964_io_out_0; // @[MUL.scala 125:16]
  assign m_2148_io_in_1 = m_1963_io_out_1; // @[MUL.scala 126:16]
  assign m_2149_io_in_0 = m_1965_io_out_0; // @[MUL.scala 125:16]
  assign m_2149_io_in_1 = m_1964_io_out_1; // @[MUL.scala 126:16]
  assign m_2150_io_in_0 = m_1966_io_out_0; // @[MUL.scala 125:16]
  assign m_2150_io_in_1 = m_1965_io_out_1; // @[MUL.scala 126:16]
  assign m_2151_io_in_0 = m_1967_io_s; // @[MUL.scala 252:21]
  assign m_2151_io_in_1 = m_1966_io_out_1; // @[MUL.scala 126:16]
  assign m_2152_io_in_0 = m_1968_io_s; // @[MUL.scala 252:21]
  assign m_2152_io_in_1 = m_1967_io_cout; // @[MUL.scala 253:22]
  assign m_2153_io_in_0 = m_1969_io_s; // @[MUL.scala 252:21]
  assign m_2153_io_in_1 = m_1968_io_cout; // @[MUL.scala 253:22]
  assign m_2154_io_in_0 = m_1970_io_s; // @[MUL.scala 252:21]
  assign m_2154_io_in_1 = m_1969_io_cout; // @[MUL.scala 253:22]
  assign m_2155_io_in_0 = m_1971_io_s; // @[MUL.scala 252:21]
  assign m_2155_io_in_1 = m_1970_io_cout; // @[MUL.scala 253:22]
  assign m_2156_io_in_0 = m_1972_io_s; // @[MUL.scala 252:21]
  assign m_2156_io_in_1 = m_1971_io_cout; // @[MUL.scala 253:22]
  assign m_2157_io_in_0 = m_1973_io_s; // @[MUL.scala 252:21]
  assign m_2157_io_in_1 = m_1972_io_cout; // @[MUL.scala 253:22]
  assign m_2158_io_in_0 = m_1974_io_s; // @[MUL.scala 252:21]
  assign m_2158_io_in_1 = m_1973_io_cout; // @[MUL.scala 253:22]
  assign m_2159_io_in_0 = m_1975_io_s; // @[MUL.scala 252:21]
  assign m_2159_io_in_1 = m_1974_io_cout; // @[MUL.scala 253:22]
  assign m_2160_io_x1 = m_1976_io_s; // @[MUL.scala 252:21]
  assign m_2160_io_x2 = m_1975_io_cout; // @[MUL.scala 253:22]
  assign m_2160_io_x3 = r_2368; // @[MUL.scala 105:13]
  assign m_2161_io_x1 = m_1977_io_s; // @[MUL.scala 252:21]
  assign m_2161_io_x2 = m_1976_io_cout; // @[MUL.scala 253:22]
  assign m_2161_io_x3 = r_2372; // @[MUL.scala 105:13]
  assign m_2162_io_x1 = m_1978_io_s; // @[MUL.scala 252:21]
  assign m_2162_io_x2 = m_1977_io_cout; // @[MUL.scala 253:22]
  assign m_2162_io_x3 = r_2376; // @[MUL.scala 105:13]
  assign m_2163_io_x1 = m_1979_io_s; // @[MUL.scala 252:21]
  assign m_2163_io_x2 = m_1978_io_cout; // @[MUL.scala 253:22]
  assign m_2163_io_x3 = r_2380; // @[MUL.scala 105:13]
  assign m_2164_io_x1 = m_1980_io_s; // @[MUL.scala 252:21]
  assign m_2164_io_x2 = m_1979_io_cout; // @[MUL.scala 253:22]
  assign m_2164_io_x3 = r_2384; // @[MUL.scala 105:13]
  assign m_2165_io_x1 = m_1981_io_s; // @[MUL.scala 252:21]
  assign m_2165_io_x2 = m_1980_io_cout; // @[MUL.scala 253:22]
  assign m_2165_io_x3 = r_2388; // @[MUL.scala 105:13]
  assign m_2166_io_x1 = m_1982_io_s; // @[MUL.scala 252:21]
  assign m_2166_io_x2 = m_1981_io_cout; // @[MUL.scala 253:22]
  assign m_2166_io_x3 = r_2392; // @[MUL.scala 105:13]
  assign m_2167_io_x1 = m_1983_io_s; // @[MUL.scala 252:21]
  assign m_2167_io_x2 = m_1982_io_cout; // @[MUL.scala 253:22]
  assign m_2167_io_x3 = r_2396; // @[MUL.scala 105:13]
  assign m_2168_io_x1 = m_1984_io_s; // @[MUL.scala 252:21]
  assign m_2168_io_x2 = m_1983_io_cout; // @[MUL.scala 253:22]
  assign m_2168_io_x3 = r_2400; // @[MUL.scala 105:13]
  assign m_2169_io_x1 = m_1985_io_s; // @[MUL.scala 252:21]
  assign m_2169_io_x2 = m_1984_io_cout; // @[MUL.scala 253:22]
  assign m_2169_io_x3 = r_2404; // @[MUL.scala 105:13]
  assign m_2170_io_x1 = m_1986_io_s; // @[MUL.scala 252:21]
  assign m_2170_io_x2 = m_1985_io_cout; // @[MUL.scala 253:22]
  assign m_2170_io_x3 = r_2408; // @[MUL.scala 105:13]
  assign m_2171_io_x1 = m_1987_io_s; // @[MUL.scala 252:21]
  assign m_2171_io_x2 = m_1986_io_cout; // @[MUL.scala 253:22]
  assign m_2171_io_x3 = r_2412; // @[MUL.scala 105:13]
  assign m_2172_io_x1 = m_1988_io_s; // @[MUL.scala 252:21]
  assign m_2172_io_x2 = m_1987_io_cout; // @[MUL.scala 253:22]
  assign m_2172_io_x3 = m_1989_io_out_0; // @[MUL.scala 105:13]
  assign m_2173_io_x1 = m_1990_io_s; // @[MUL.scala 252:21]
  assign m_2173_io_x2 = m_1988_io_cout; // @[MUL.scala 253:22]
  assign m_2173_io_x3 = m_1991_io_out_0; // @[MUL.scala 105:13]
  assign m_2174_io_x1 = m_1992_io_s; // @[MUL.scala 252:21]
  assign m_2174_io_x2 = m_1990_io_cout; // @[MUL.scala 253:22]
  assign m_2174_io_x3 = m_1993_io_out_0; // @[MUL.scala 105:13]
  assign m_2175_io_x1 = m_1994_io_s; // @[MUL.scala 252:21]
  assign m_2175_io_x2 = m_1992_io_cout; // @[MUL.scala 253:22]
  assign m_2175_io_x3 = m_1995_io_out_0; // @[MUL.scala 105:13]
  assign m_2176_io_x1 = m_1996_io_s; // @[MUL.scala 252:21]
  assign m_2176_io_x2 = m_1994_io_cout; // @[MUL.scala 253:22]
  assign m_2176_io_x3 = m_1997_io_out_0; // @[MUL.scala 105:13]
  assign m_2177_io_x1 = m_1998_io_s; // @[MUL.scala 252:21]
  assign m_2177_io_x2 = m_1996_io_cout; // @[MUL.scala 253:22]
  assign m_2177_io_x3 = m_1999_io_out_0; // @[MUL.scala 105:13]
  assign m_2178_io_x1 = m_2000_io_s; // @[MUL.scala 252:21]
  assign m_2178_io_x2 = m_1998_io_cout; // @[MUL.scala 253:22]
  assign m_2178_io_x3 = m_2001_io_out_0; // @[MUL.scala 105:13]
  assign m_2179_io_x1 = m_2002_io_s; // @[MUL.scala 252:21]
  assign m_2179_io_x2 = m_2000_io_cout; // @[MUL.scala 253:22]
  assign m_2179_io_x3 = m_2003_io_s; // @[MUL.scala 252:21]
  assign m_2180_io_x1 = m_2004_io_s; // @[MUL.scala 252:21]
  assign m_2180_io_x2 = m_2002_io_cout; // @[MUL.scala 253:22]
  assign m_2180_io_x3 = m_2005_io_s; // @[MUL.scala 252:21]
  assign m_2181_io_x1 = m_2006_io_s; // @[MUL.scala 252:21]
  assign m_2181_io_x2 = m_2004_io_cout; // @[MUL.scala 253:22]
  assign m_2181_io_x3 = m_2007_io_s; // @[MUL.scala 252:21]
  assign m_2182_io_x1 = m_2008_io_s; // @[MUL.scala 252:21]
  assign m_2182_io_x2 = m_2006_io_cout; // @[MUL.scala 253:22]
  assign m_2182_io_x3 = m_2009_io_s; // @[MUL.scala 252:21]
  assign m_2183_io_x1 = m_2010_io_s; // @[MUL.scala 252:21]
  assign m_2183_io_x2 = m_2008_io_cout; // @[MUL.scala 253:22]
  assign m_2183_io_x3 = m_2011_io_s; // @[MUL.scala 252:21]
  assign m_2184_io_x1 = m_2012_io_s; // @[MUL.scala 252:21]
  assign m_2184_io_x2 = m_2010_io_cout; // @[MUL.scala 253:22]
  assign m_2184_io_x3 = m_2013_io_s; // @[MUL.scala 252:21]
  assign m_2185_io_x1 = m_2014_io_s; // @[MUL.scala 252:21]
  assign m_2185_io_x2 = m_2012_io_cout; // @[MUL.scala 253:22]
  assign m_2185_io_x3 = m_2015_io_s; // @[MUL.scala 252:21]
  assign m_2186_io_x1 = m_2016_io_s; // @[MUL.scala 252:21]
  assign m_2186_io_x2 = m_2014_io_cout; // @[MUL.scala 253:22]
  assign m_2186_io_x3 = m_2017_io_s; // @[MUL.scala 252:21]
  assign m_2187_io_x1 = m_2018_io_s; // @[MUL.scala 252:21]
  assign m_2187_io_x2 = m_2016_io_cout; // @[MUL.scala 253:22]
  assign m_2187_io_x3 = m_2019_io_s; // @[MUL.scala 252:21]
  assign m_2188_io_x1 = m_2020_io_s; // @[MUL.scala 252:21]
  assign m_2188_io_x2 = m_2018_io_cout; // @[MUL.scala 253:22]
  assign m_2188_io_x3 = m_2021_io_s; // @[MUL.scala 252:21]
  assign m_2189_io_x1 = m_2022_io_s; // @[MUL.scala 252:21]
  assign m_2189_io_x2 = m_2020_io_cout; // @[MUL.scala 253:22]
  assign m_2189_io_x3 = m_2023_io_s; // @[MUL.scala 252:21]
  assign m_2190_io_x1 = m_2024_io_s; // @[MUL.scala 252:21]
  assign m_2190_io_x2 = m_2022_io_cout; // @[MUL.scala 253:22]
  assign m_2190_io_x3 = m_2025_io_s; // @[MUL.scala 252:21]
  assign m_2191_io_x1 = m_2026_io_s; // @[MUL.scala 252:21]
  assign m_2191_io_x2 = m_2024_io_cout; // @[MUL.scala 253:22]
  assign m_2191_io_x3 = m_2027_io_s; // @[MUL.scala 252:21]
  assign m_2192_io_in_0 = m_2025_io_cout; // @[MUL.scala 253:22]
  assign m_2192_io_in_1 = r_2526; // @[MUL.scala 126:16]
  assign m_2193_io_x1 = m_2028_io_s; // @[MUL.scala 252:21]
  assign m_2193_io_x2 = m_2026_io_cout; // @[MUL.scala 253:22]
  assign m_2193_io_x3 = m_2029_io_s; // @[MUL.scala 252:21]
  assign m_2194_io_in_0 = m_2027_io_cout; // @[MUL.scala 253:22]
  assign m_2194_io_in_1 = r_2533; // @[MUL.scala 126:16]
  assign m_2195_io_x1 = m_2030_io_s; // @[MUL.scala 252:21]
  assign m_2195_io_x2 = m_2028_io_cout; // @[MUL.scala 253:22]
  assign m_2195_io_x3 = m_2031_io_s; // @[MUL.scala 252:21]
  assign m_2196_io_in_0 = m_2029_io_cout; // @[MUL.scala 253:22]
  assign m_2196_io_in_1 = r_2540; // @[MUL.scala 126:16]
  assign m_2197_io_x1 = m_2032_io_s; // @[MUL.scala 252:21]
  assign m_2197_io_x2 = m_2030_io_cout; // @[MUL.scala 253:22]
  assign m_2197_io_x3 = m_2033_io_s; // @[MUL.scala 252:21]
  assign m_2198_io_in_0 = m_2031_io_cout; // @[MUL.scala 253:22]
  assign m_2198_io_in_1 = r_2547; // @[MUL.scala 126:16]
  assign m_2199_io_x1 = m_2034_io_s; // @[MUL.scala 252:21]
  assign m_2199_io_x2 = m_2032_io_cout; // @[MUL.scala 253:22]
  assign m_2199_io_x3 = m_2035_io_s; // @[MUL.scala 252:21]
  assign m_2200_io_in_0 = m_2033_io_cout; // @[MUL.scala 253:22]
  assign m_2200_io_in_1 = r_2554; // @[MUL.scala 126:16]
  assign m_2201_io_x1 = m_2036_io_s; // @[MUL.scala 252:21]
  assign m_2201_io_x2 = m_2034_io_cout; // @[MUL.scala 253:22]
  assign m_2201_io_x3 = m_2037_io_s; // @[MUL.scala 252:21]
  assign m_2202_io_in_0 = m_2035_io_cout; // @[MUL.scala 253:22]
  assign m_2202_io_in_1 = r_2561; // @[MUL.scala 126:16]
  assign m_2203_io_x1 = m_2038_io_s; // @[MUL.scala 252:21]
  assign m_2203_io_x2 = m_2036_io_cout; // @[MUL.scala 253:22]
  assign m_2203_io_x3 = m_2039_io_s; // @[MUL.scala 252:21]
  assign m_2204_io_in_0 = m_2037_io_cout; // @[MUL.scala 253:22]
  assign m_2204_io_in_1 = r_2568; // @[MUL.scala 126:16]
  assign m_2205_io_x1 = m_2040_io_s; // @[MUL.scala 252:21]
  assign m_2205_io_x2 = m_2038_io_cout; // @[MUL.scala 253:22]
  assign m_2205_io_x3 = m_2041_io_s; // @[MUL.scala 252:21]
  assign m_2206_io_in_0 = m_2039_io_cout; // @[MUL.scala 253:22]
  assign m_2206_io_in_1 = r_2575; // @[MUL.scala 126:16]
  assign m_2207_io_x1 = m_2042_io_s; // @[MUL.scala 252:21]
  assign m_2207_io_x2 = m_2040_io_cout; // @[MUL.scala 253:22]
  assign m_2207_io_x3 = m_2043_io_s; // @[MUL.scala 252:21]
  assign m_2208_io_in_0 = m_2041_io_cout; // @[MUL.scala 253:22]
  assign m_2208_io_in_1 = r_2582; // @[MUL.scala 126:16]
  assign m_2209_io_x1 = m_2044_io_s; // @[MUL.scala 252:21]
  assign m_2209_io_x2 = m_2042_io_cout; // @[MUL.scala 253:22]
  assign m_2209_io_x3 = m_2045_io_s; // @[MUL.scala 252:21]
  assign m_2210_io_in_0 = m_2043_io_cout; // @[MUL.scala 253:22]
  assign m_2210_io_in_1 = r_2589; // @[MUL.scala 126:16]
  assign m_2211_io_x1 = m_2046_io_s; // @[MUL.scala 252:21]
  assign m_2211_io_x2 = m_2044_io_cout; // @[MUL.scala 253:22]
  assign m_2211_io_x3 = m_2047_io_s; // @[MUL.scala 252:21]
  assign m_2212_io_in_0 = m_2045_io_cout; // @[MUL.scala 253:22]
  assign m_2212_io_in_1 = r_2596; // @[MUL.scala 126:16]
  assign m_2213_io_x1 = m_2048_io_s; // @[MUL.scala 252:21]
  assign m_2213_io_x2 = m_2046_io_cout; // @[MUL.scala 253:22]
  assign m_2213_io_x3 = m_2049_io_s; // @[MUL.scala 252:21]
  assign m_2214_io_in_0 = m_2047_io_cout; // @[MUL.scala 253:22]
  assign m_2214_io_in_1 = r_2603; // @[MUL.scala 126:16]
  assign m_2215_io_x1 = m_2050_io_s; // @[MUL.scala 252:21]
  assign m_2215_io_x2 = m_2048_io_cout; // @[MUL.scala 253:22]
  assign m_2215_io_x3 = m_2051_io_s; // @[MUL.scala 252:21]
  assign m_2216_io_in_0 = m_2049_io_cout; // @[MUL.scala 253:22]
  assign m_2216_io_in_1 = r_2610; // @[MUL.scala 126:16]
  assign m_2217_io_x1 = m_2052_io_s; // @[MUL.scala 252:21]
  assign m_2217_io_x2 = m_2050_io_cout; // @[MUL.scala 253:22]
  assign m_2217_io_x3 = m_2053_io_s; // @[MUL.scala 252:21]
  assign m_2218_io_in_0 = m_2051_io_cout; // @[MUL.scala 253:22]
  assign m_2218_io_in_1 = r_2617; // @[MUL.scala 126:16]
  assign m_2219_io_x1 = m_2054_io_s; // @[MUL.scala 252:21]
  assign m_2219_io_x2 = m_2052_io_cout; // @[MUL.scala 253:22]
  assign m_2219_io_x3 = m_2055_io_s; // @[MUL.scala 252:21]
  assign m_2220_io_in_0 = m_2053_io_cout; // @[MUL.scala 253:22]
  assign m_2220_io_in_1 = r_2624; // @[MUL.scala 126:16]
  assign m_2221_io_x1 = m_2056_io_s; // @[MUL.scala 252:21]
  assign m_2221_io_x2 = m_2054_io_cout; // @[MUL.scala 253:22]
  assign m_2221_io_x3 = m_2057_io_s; // @[MUL.scala 252:21]
  assign m_2222_io_in_0 = m_2055_io_cout; // @[MUL.scala 253:22]
  assign m_2222_io_in_1 = r_2631; // @[MUL.scala 126:16]
  assign m_2223_io_x1 = m_2058_io_s; // @[MUL.scala 252:21]
  assign m_2223_io_x2 = m_2056_io_cout; // @[MUL.scala 253:22]
  assign m_2223_io_x3 = m_2059_io_s; // @[MUL.scala 252:21]
  assign m_2224_io_in_0 = m_2057_io_cout; // @[MUL.scala 253:22]
  assign m_2224_io_in_1 = r_2638; // @[MUL.scala 126:16]
  assign m_2225_io_x1 = m_2060_io_s; // @[MUL.scala 252:21]
  assign m_2225_io_x2 = m_2058_io_cout; // @[MUL.scala 253:22]
  assign m_2225_io_x3 = m_2061_io_s; // @[MUL.scala 252:21]
  assign m_2226_io_in_0 = m_2059_io_cout; // @[MUL.scala 253:22]
  assign m_2226_io_in_1 = r_2645; // @[MUL.scala 126:16]
  assign m_2227_io_x1 = m_2062_io_s; // @[MUL.scala 252:21]
  assign m_2227_io_x2 = m_2060_io_cout; // @[MUL.scala 253:22]
  assign m_2227_io_x3 = m_2063_io_s; // @[MUL.scala 252:21]
  assign m_2228_io_in_0 = m_2061_io_cout; // @[MUL.scala 253:22]
  assign m_2228_io_in_1 = r_2652; // @[MUL.scala 126:16]
  assign m_2229_io_x1 = m_2064_io_s; // @[MUL.scala 252:21]
  assign m_2229_io_x2 = m_2062_io_cout; // @[MUL.scala 253:22]
  assign m_2229_io_x3 = m_2065_io_s; // @[MUL.scala 252:21]
  assign m_2230_io_in_0 = m_2063_io_cout; // @[MUL.scala 253:22]
  assign m_2230_io_in_1 = r_2659; // @[MUL.scala 126:16]
  assign m_2231_io_x1 = m_2066_io_s; // @[MUL.scala 252:21]
  assign m_2231_io_x2 = m_2064_io_cout; // @[MUL.scala 253:22]
  assign m_2231_io_x3 = m_2067_io_s; // @[MUL.scala 252:21]
  assign m_2232_io_in_0 = m_2065_io_cout; // @[MUL.scala 253:22]
  assign m_2232_io_in_1 = r_2666; // @[MUL.scala 126:16]
  assign m_2233_io_x1 = m_2068_io_s; // @[MUL.scala 252:21]
  assign m_2233_io_x2 = m_2066_io_cout; // @[MUL.scala 253:22]
  assign m_2233_io_x3 = m_2069_io_s; // @[MUL.scala 252:21]
  assign m_2234_io_x1 = m_2070_io_s; // @[MUL.scala 252:21]
  assign m_2234_io_x2 = m_2068_io_cout; // @[MUL.scala 253:22]
  assign m_2234_io_x3 = m_2071_io_s; // @[MUL.scala 252:21]
  assign m_2235_io_x1 = m_2072_io_s; // @[MUL.scala 252:21]
  assign m_2235_io_x2 = m_2070_io_cout; // @[MUL.scala 253:22]
  assign m_2235_io_x3 = m_2073_io_s; // @[MUL.scala 252:21]
  assign m_2236_io_x1 = m_2074_io_s; // @[MUL.scala 252:21]
  assign m_2236_io_x2 = m_2072_io_cout; // @[MUL.scala 253:22]
  assign m_2236_io_x3 = m_2075_io_s; // @[MUL.scala 252:21]
  assign m_2237_io_x1 = m_2076_io_s; // @[MUL.scala 252:21]
  assign m_2237_io_x2 = m_2074_io_cout; // @[MUL.scala 253:22]
  assign m_2237_io_x3 = m_2077_io_s; // @[MUL.scala 252:21]
  assign m_2238_io_x1 = m_2078_io_s; // @[MUL.scala 252:21]
  assign m_2238_io_x2 = m_2076_io_cout; // @[MUL.scala 253:22]
  assign m_2238_io_x3 = m_2079_io_s; // @[MUL.scala 252:21]
  assign m_2239_io_x1 = m_2080_io_s; // @[MUL.scala 252:21]
  assign m_2239_io_x2 = m_2078_io_cout; // @[MUL.scala 253:22]
  assign m_2239_io_x3 = m_2081_io_s; // @[MUL.scala 252:21]
  assign m_2240_io_x1 = m_2082_io_s; // @[MUL.scala 252:21]
  assign m_2240_io_x2 = m_2080_io_cout; // @[MUL.scala 253:22]
  assign m_2240_io_x3 = m_2083_io_s; // @[MUL.scala 252:21]
  assign m_2241_io_x1 = m_2084_io_s; // @[MUL.scala 252:21]
  assign m_2241_io_x2 = m_2082_io_cout; // @[MUL.scala 253:22]
  assign m_2241_io_x3 = m_2085_io_s; // @[MUL.scala 252:21]
  assign m_2242_io_x1 = m_2086_io_s; // @[MUL.scala 252:21]
  assign m_2242_io_x2 = m_2084_io_cout; // @[MUL.scala 253:22]
  assign m_2242_io_x3 = m_2087_io_s; // @[MUL.scala 252:21]
  assign m_2243_io_x1 = m_2088_io_s; // @[MUL.scala 252:21]
  assign m_2243_io_x2 = m_2086_io_cout; // @[MUL.scala 253:22]
  assign m_2243_io_x3 = m_2089_io_s; // @[MUL.scala 252:21]
  assign m_2244_io_x1 = m_2090_io_s; // @[MUL.scala 252:21]
  assign m_2244_io_x2 = m_2088_io_cout; // @[MUL.scala 253:22]
  assign m_2244_io_x3 = m_2091_io_s; // @[MUL.scala 252:21]
  assign m_2245_io_x1 = m_2092_io_s; // @[MUL.scala 252:21]
  assign m_2245_io_x2 = m_2090_io_cout; // @[MUL.scala 253:22]
  assign m_2245_io_x3 = m_2093_io_s; // @[MUL.scala 252:21]
  assign m_2246_io_x1 = m_2094_io_s; // @[MUL.scala 252:21]
  assign m_2246_io_x2 = m_2092_io_cout; // @[MUL.scala 253:22]
  assign m_2246_io_x3 = m_2095_io_out_0; // @[MUL.scala 105:13]
  assign m_2247_io_x1 = m_2096_io_s; // @[MUL.scala 252:21]
  assign m_2247_io_x2 = m_2094_io_cout; // @[MUL.scala 253:22]
  assign m_2247_io_x3 = m_2097_io_out_0; // @[MUL.scala 105:13]
  assign m_2248_io_x1 = m_2098_io_s; // @[MUL.scala 252:21]
  assign m_2248_io_x2 = m_2096_io_cout; // @[MUL.scala 253:22]
  assign m_2248_io_x3 = m_2099_io_out_0; // @[MUL.scala 105:13]
  assign m_2249_io_x1 = m_2100_io_s; // @[MUL.scala 252:21]
  assign m_2249_io_x2 = m_2098_io_cout; // @[MUL.scala 253:22]
  assign m_2249_io_x3 = m_2101_io_out_0; // @[MUL.scala 105:13]
  assign m_2250_io_x1 = m_2102_io_s; // @[MUL.scala 252:21]
  assign m_2250_io_x2 = m_2100_io_cout; // @[MUL.scala 253:22]
  assign m_2250_io_x3 = m_2103_io_out_0; // @[MUL.scala 105:13]
  assign m_2251_io_x1 = m_2104_io_s; // @[MUL.scala 252:21]
  assign m_2251_io_x2 = m_2102_io_cout; // @[MUL.scala 253:22]
  assign m_2251_io_x3 = r_2773; // @[MUL.scala 105:13]
  assign m_2252_io_x1 = m_2105_io_s; // @[MUL.scala 252:21]
  assign m_2252_io_x2 = m_2104_io_cout; // @[MUL.scala 253:22]
  assign m_2252_io_x3 = r_2777; // @[MUL.scala 105:13]
  assign m_2253_io_x1 = m_2106_io_s; // @[MUL.scala 252:21]
  assign m_2253_io_x2 = m_2105_io_cout; // @[MUL.scala 253:22]
  assign m_2253_io_x3 = r_2781; // @[MUL.scala 105:13]
  assign m_2254_io_x1 = m_2107_io_s; // @[MUL.scala 252:21]
  assign m_2254_io_x2 = m_2106_io_cout; // @[MUL.scala 253:22]
  assign m_2254_io_x3 = r_2785; // @[MUL.scala 105:13]
  assign m_2255_io_x1 = m_2108_io_s; // @[MUL.scala 252:21]
  assign m_2255_io_x2 = m_2107_io_cout; // @[MUL.scala 253:22]
  assign m_2255_io_x3 = r_2789; // @[MUL.scala 105:13]
  assign m_2256_io_x1 = m_2109_io_s; // @[MUL.scala 252:21]
  assign m_2256_io_x2 = m_2108_io_cout; // @[MUL.scala 253:22]
  assign m_2256_io_x3 = r_2793; // @[MUL.scala 105:13]
  assign m_2257_io_x1 = m_2110_io_s; // @[MUL.scala 252:21]
  assign m_2257_io_x2 = m_2109_io_cout; // @[MUL.scala 253:22]
  assign m_2257_io_x3 = r_2797; // @[MUL.scala 105:13]
  assign m_2258_io_x1 = m_2111_io_s; // @[MUL.scala 252:21]
  assign m_2258_io_x2 = m_2110_io_cout; // @[MUL.scala 253:22]
  assign m_2258_io_x3 = r_2801; // @[MUL.scala 105:13]
  assign m_2259_io_x1 = m_2112_io_s; // @[MUL.scala 252:21]
  assign m_2259_io_x2 = m_2111_io_cout; // @[MUL.scala 253:22]
  assign m_2259_io_x3 = r_2805; // @[MUL.scala 105:13]
  assign m_2260_io_x1 = m_2113_io_s; // @[MUL.scala 252:21]
  assign m_2260_io_x2 = m_2112_io_cout; // @[MUL.scala 253:22]
  assign m_2260_io_x3 = r_2809; // @[MUL.scala 105:13]
  assign m_2261_io_x1 = m_2114_io_s; // @[MUL.scala 252:21]
  assign m_2261_io_x2 = m_2113_io_cout; // @[MUL.scala 253:22]
  assign m_2261_io_x3 = r_2813; // @[MUL.scala 105:13]
  assign m_2262_io_x1 = m_2115_io_s; // @[MUL.scala 252:21]
  assign m_2262_io_x2 = m_2114_io_cout; // @[MUL.scala 253:22]
  assign m_2262_io_x3 = r_2817; // @[MUL.scala 105:13]
  assign m_2263_io_in_0 = m_2116_io_s; // @[MUL.scala 252:21]
  assign m_2263_io_in_1 = m_2115_io_cout; // @[MUL.scala 253:22]
  assign m_2264_io_in_0 = m_2117_io_s; // @[MUL.scala 252:21]
  assign m_2264_io_in_1 = m_2116_io_cout; // @[MUL.scala 253:22]
  assign m_2265_io_in_0 = m_2118_io_s; // @[MUL.scala 252:21]
  assign m_2265_io_in_1 = m_2117_io_cout; // @[MUL.scala 253:22]
  assign m_2266_io_in_0 = m_2119_io_s; // @[MUL.scala 252:21]
  assign m_2266_io_in_1 = m_2118_io_cout; // @[MUL.scala 253:22]
  assign m_2267_io_in_0 = m_2120_io_s; // @[MUL.scala 252:21]
  assign m_2267_io_in_1 = m_2119_io_cout; // @[MUL.scala 253:22]
  assign m_2268_io_in_0 = m_2121_io_s; // @[MUL.scala 252:21]
  assign m_2268_io_in_1 = m_2120_io_cout; // @[MUL.scala 253:22]
  assign m_2269_io_in_0 = m_2122_io_s; // @[MUL.scala 252:21]
  assign m_2269_io_in_1 = m_2121_io_cout; // @[MUL.scala 253:22]
  assign m_2270_io_in_0 = m_2123_io_out_0; // @[MUL.scala 125:16]
  assign m_2270_io_in_1 = m_2122_io_cout; // @[MUL.scala 253:22]
  assign m_2271_io_in_0 = m_2124_io_out_0; // @[MUL.scala 125:16]
  assign m_2271_io_in_1 = m_2123_io_out_1; // @[MUL.scala 126:16]
  assign m_2272_io_in_0 = m_2125_io_out_0; // @[MUL.scala 125:16]
  assign m_2272_io_in_1 = m_2124_io_out_1; // @[MUL.scala 126:16]
  assign m_2273_io_in_0 = m_2126_io_out_0; // @[MUL.scala 125:16]
  assign m_2273_io_in_1 = m_2125_io_out_1; // @[MUL.scala 126:16]
  assign m_2274_io_in_0 = m_2127_io_out_0; // @[MUL.scala 125:16]
  assign m_2274_io_in_1 = m_2126_io_out_1; // @[MUL.scala 126:16]
  assign m_2275_io_in_0 = m_2128_io_out_0; // @[MUL.scala 125:16]
  assign m_2275_io_in_1 = m_2127_io_out_1; // @[MUL.scala 126:16]
  assign m_2276_io_in_0 = m_2129_io_out_0; // @[MUL.scala 125:16]
  assign m_2276_io_in_1 = m_2128_io_out_1; // @[MUL.scala 126:16]
  assign m_2277_io_in_0 = m_2130_io_out_0; // @[MUL.scala 125:16]
  assign m_2277_io_in_1 = m_2129_io_out_1; // @[MUL.scala 126:16]
  assign m_2278_io_in_0 = m_2131_io_out_0; // @[MUL.scala 125:16]
  assign m_2278_io_in_1 = m_2130_io_out_1; // @[MUL.scala 126:16]
  assign m_2279_io_in_0 = m_2132_io_out_0; // @[MUL.scala 125:16]
  assign m_2279_io_in_1 = m_2131_io_out_1; // @[MUL.scala 126:16]
  assign m_2280_io_in_0 = m_2133_io_out_0; // @[MUL.scala 125:16]
  assign m_2280_io_in_1 = m_2132_io_out_1; // @[MUL.scala 126:16]
  assign m_2281_io_in_0 = m_2134_io_out_0; // @[MUL.scala 125:16]
  assign m_2281_io_in_1 = m_2133_io_out_1; // @[MUL.scala 126:16]
  assign m_2282_io_in_0 = m_2135_io_out_0; // @[MUL.scala 125:16]
  assign m_2282_io_in_1 = m_2134_io_out_1; // @[MUL.scala 126:16]
  assign m_2283_io_in_0 = m_2136_io_out_0; // @[MUL.scala 125:16]
  assign m_2283_io_in_1 = m_2135_io_out_1; // @[MUL.scala 126:16]
  assign m_2284_io_in_0 = m_2137_io_out_0; // @[MUL.scala 125:16]
  assign m_2284_io_in_1 = m_2136_io_out_1; // @[MUL.scala 126:16]
  assign m_2285_io_in_0 = m_2138_io_out_0; // @[MUL.scala 125:16]
  assign m_2285_io_in_1 = m_2137_io_out_1; // @[MUL.scala 126:16]
  assign m_2286_io_in_0 = m_2140_io_out_0; // @[MUL.scala 125:16]
  assign m_2286_io_in_1 = m_2139_io_out_1; // @[MUL.scala 126:16]
  assign m_2287_io_in_0 = m_2141_io_out_0; // @[MUL.scala 125:16]
  assign m_2287_io_in_1 = m_2140_io_out_1; // @[MUL.scala 126:16]
  assign m_2288_io_in_0 = m_2142_io_out_0; // @[MUL.scala 125:16]
  assign m_2288_io_in_1 = m_2141_io_out_1; // @[MUL.scala 126:16]
  assign m_2289_io_in_0 = m_2143_io_out_0; // @[MUL.scala 125:16]
  assign m_2289_io_in_1 = m_2142_io_out_1; // @[MUL.scala 126:16]
  assign m_2290_io_in_0 = m_2144_io_out_0; // @[MUL.scala 125:16]
  assign m_2290_io_in_1 = m_2143_io_out_1; // @[MUL.scala 126:16]
  assign m_2291_io_in_0 = m_2145_io_out_0; // @[MUL.scala 125:16]
  assign m_2291_io_in_1 = m_2144_io_out_1; // @[MUL.scala 126:16]
  assign m_2292_io_in_0 = m_2146_io_out_0; // @[MUL.scala 125:16]
  assign m_2292_io_in_1 = m_2145_io_out_1; // @[MUL.scala 126:16]
  assign m_2293_io_in_0 = m_2147_io_out_0; // @[MUL.scala 125:16]
  assign m_2293_io_in_1 = m_2146_io_out_1; // @[MUL.scala 126:16]
  assign m_2294_io_in_0 = m_2148_io_out_0; // @[MUL.scala 125:16]
  assign m_2294_io_in_1 = m_2147_io_out_1; // @[MUL.scala 126:16]
  assign m_2295_io_in_0 = m_2149_io_out_0; // @[MUL.scala 125:16]
  assign m_2295_io_in_1 = m_2148_io_out_1; // @[MUL.scala 126:16]
  assign m_2296_io_in_0 = m_2150_io_out_0; // @[MUL.scala 125:16]
  assign m_2296_io_in_1 = m_2149_io_out_1; // @[MUL.scala 126:16]
  assign m_2297_io_in_0 = m_2151_io_out_0; // @[MUL.scala 125:16]
  assign m_2297_io_in_1 = m_2150_io_out_1; // @[MUL.scala 126:16]
  assign m_2298_io_in_0 = m_2152_io_out_0; // @[MUL.scala 125:16]
  assign m_2298_io_in_1 = m_2151_io_out_1; // @[MUL.scala 126:16]
  assign m_2299_io_in_0 = m_2153_io_out_0; // @[MUL.scala 125:16]
  assign m_2299_io_in_1 = m_2152_io_out_1; // @[MUL.scala 126:16]
  assign m_2300_io_in_0 = m_2154_io_out_0; // @[MUL.scala 125:16]
  assign m_2300_io_in_1 = m_2153_io_out_1; // @[MUL.scala 126:16]
  assign m_2301_io_in_0 = m_2155_io_out_0; // @[MUL.scala 125:16]
  assign m_2301_io_in_1 = m_2154_io_out_1; // @[MUL.scala 126:16]
  assign m_2302_io_in_0 = m_2156_io_out_0; // @[MUL.scala 125:16]
  assign m_2302_io_in_1 = m_2155_io_out_1; // @[MUL.scala 126:16]
  assign m_2303_io_in_0 = m_2157_io_out_0; // @[MUL.scala 125:16]
  assign m_2303_io_in_1 = m_2156_io_out_1; // @[MUL.scala 126:16]
  assign m_2304_io_in_0 = m_2158_io_out_0; // @[MUL.scala 125:16]
  assign m_2304_io_in_1 = m_2157_io_out_1; // @[MUL.scala 126:16]
  assign m_2305_io_in_0 = m_2159_io_out_0; // @[MUL.scala 125:16]
  assign m_2305_io_in_1 = m_2158_io_out_1; // @[MUL.scala 126:16]
  assign m_2306_io_in_0 = m_2160_io_s; // @[MUL.scala 252:21]
  assign m_2306_io_in_1 = m_2159_io_out_1; // @[MUL.scala 126:16]
  assign m_2307_io_in_0 = m_2161_io_s; // @[MUL.scala 252:21]
  assign m_2307_io_in_1 = m_2160_io_cout; // @[MUL.scala 253:22]
  assign m_2308_io_in_0 = m_2162_io_s; // @[MUL.scala 252:21]
  assign m_2308_io_in_1 = m_2161_io_cout; // @[MUL.scala 253:22]
  assign m_2309_io_in_0 = m_2163_io_s; // @[MUL.scala 252:21]
  assign m_2309_io_in_1 = m_2162_io_cout; // @[MUL.scala 253:22]
  assign m_2310_io_in_0 = m_2164_io_s; // @[MUL.scala 252:21]
  assign m_2310_io_in_1 = m_2163_io_cout; // @[MUL.scala 253:22]
  assign m_2311_io_in_0 = m_2165_io_s; // @[MUL.scala 252:21]
  assign m_2311_io_in_1 = m_2164_io_cout; // @[MUL.scala 253:22]
  assign m_2312_io_in_0 = m_2166_io_s; // @[MUL.scala 252:21]
  assign m_2312_io_in_1 = m_2165_io_cout; // @[MUL.scala 253:22]
  assign m_2313_io_in_0 = m_2167_io_s; // @[MUL.scala 252:21]
  assign m_2313_io_in_1 = m_2166_io_cout; // @[MUL.scala 253:22]
  assign m_2314_io_in_0 = m_2168_io_s; // @[MUL.scala 252:21]
  assign m_2314_io_in_1 = m_2167_io_cout; // @[MUL.scala 253:22]
  assign m_2315_io_in_0 = m_2169_io_s; // @[MUL.scala 252:21]
  assign m_2315_io_in_1 = m_2168_io_cout; // @[MUL.scala 253:22]
  assign m_2316_io_in_0 = m_2170_io_s; // @[MUL.scala 252:21]
  assign m_2316_io_in_1 = m_2169_io_cout; // @[MUL.scala 253:22]
  assign m_2317_io_in_0 = m_2171_io_s; // @[MUL.scala 252:21]
  assign m_2317_io_in_1 = m_2170_io_cout; // @[MUL.scala 253:22]
  assign m_2318_io_in_0 = m_2172_io_s; // @[MUL.scala 252:21]
  assign m_2318_io_in_1 = m_2171_io_cout; // @[MUL.scala 253:22]
  assign m_2319_io_x1 = m_2173_io_s; // @[MUL.scala 252:21]
  assign m_2319_io_x2 = m_2172_io_cout; // @[MUL.scala 253:22]
  assign m_2319_io_x3 = m_1989_io_out_1; // @[MUL.scala 105:13]
  assign m_2320_io_x1 = m_2174_io_s; // @[MUL.scala 252:21]
  assign m_2320_io_x2 = m_2173_io_cout; // @[MUL.scala 253:22]
  assign m_2320_io_x3 = m_1991_io_out_1; // @[MUL.scala 105:13]
  assign m_2321_io_x1 = m_2175_io_s; // @[MUL.scala 252:21]
  assign m_2321_io_x2 = m_2174_io_cout; // @[MUL.scala 253:22]
  assign m_2321_io_x3 = m_1993_io_out_1; // @[MUL.scala 105:13]
  assign m_2322_io_x1 = m_2176_io_s; // @[MUL.scala 252:21]
  assign m_2322_io_x2 = m_2175_io_cout; // @[MUL.scala 253:22]
  assign m_2322_io_x3 = m_1995_io_out_1; // @[MUL.scala 105:13]
  assign m_2323_io_x1 = m_2177_io_s; // @[MUL.scala 252:21]
  assign m_2323_io_x2 = m_2176_io_cout; // @[MUL.scala 253:22]
  assign m_2323_io_x3 = m_1997_io_out_1; // @[MUL.scala 105:13]
  assign m_2324_io_x1 = m_2178_io_s; // @[MUL.scala 252:21]
  assign m_2324_io_x2 = m_2177_io_cout; // @[MUL.scala 253:22]
  assign m_2324_io_x3 = m_1999_io_out_1; // @[MUL.scala 105:13]
  assign m_2325_io_x1 = m_2179_io_s; // @[MUL.scala 252:21]
  assign m_2325_io_x2 = m_2178_io_cout; // @[MUL.scala 253:22]
  assign m_2325_io_x3 = m_2001_io_out_1; // @[MUL.scala 105:13]
  assign m_2326_io_x1 = m_2180_io_s; // @[MUL.scala 252:21]
  assign m_2326_io_x2 = m_2179_io_cout; // @[MUL.scala 253:22]
  assign m_2326_io_x3 = m_2003_io_cout; // @[MUL.scala 253:22]
  assign m_2327_io_x1 = m_2181_io_s; // @[MUL.scala 252:21]
  assign m_2327_io_x2 = m_2180_io_cout; // @[MUL.scala 253:22]
  assign m_2327_io_x3 = m_2005_io_cout; // @[MUL.scala 253:22]
  assign m_2328_io_x1 = m_2182_io_s; // @[MUL.scala 252:21]
  assign m_2328_io_x2 = m_2181_io_cout; // @[MUL.scala 253:22]
  assign m_2328_io_x3 = m_2007_io_cout; // @[MUL.scala 253:22]
  assign m_2329_io_x1 = m_2183_io_s; // @[MUL.scala 252:21]
  assign m_2329_io_x2 = m_2182_io_cout; // @[MUL.scala 253:22]
  assign m_2329_io_x3 = m_2009_io_cout; // @[MUL.scala 253:22]
  assign m_2330_io_x1 = m_2184_io_s; // @[MUL.scala 252:21]
  assign m_2330_io_x2 = m_2183_io_cout; // @[MUL.scala 253:22]
  assign m_2330_io_x3 = m_2011_io_cout; // @[MUL.scala 253:22]
  assign m_2331_io_x1 = m_2185_io_s; // @[MUL.scala 252:21]
  assign m_2331_io_x2 = m_2184_io_cout; // @[MUL.scala 253:22]
  assign m_2331_io_x3 = m_2013_io_cout; // @[MUL.scala 253:22]
  assign m_2332_io_x1 = m_2186_io_s; // @[MUL.scala 252:21]
  assign m_2332_io_x2 = m_2185_io_cout; // @[MUL.scala 253:22]
  assign m_2332_io_x3 = m_2015_io_cout; // @[MUL.scala 253:22]
  assign m_2333_io_x1 = m_2187_io_s; // @[MUL.scala 252:21]
  assign m_2333_io_x2 = m_2186_io_cout; // @[MUL.scala 253:22]
  assign m_2333_io_x3 = m_2017_io_cout; // @[MUL.scala 253:22]
  assign m_2334_io_x1 = m_2188_io_s; // @[MUL.scala 252:21]
  assign m_2334_io_x2 = m_2187_io_cout; // @[MUL.scala 253:22]
  assign m_2334_io_x3 = m_2019_io_cout; // @[MUL.scala 253:22]
  assign m_2335_io_x1 = m_2189_io_s; // @[MUL.scala 252:21]
  assign m_2335_io_x2 = m_2188_io_cout; // @[MUL.scala 253:22]
  assign m_2335_io_x3 = m_2021_io_cout; // @[MUL.scala 253:22]
  assign m_2336_io_x1 = m_2190_io_s; // @[MUL.scala 252:21]
  assign m_2336_io_x2 = m_2189_io_cout; // @[MUL.scala 253:22]
  assign m_2336_io_x3 = m_2023_io_cout; // @[MUL.scala 253:22]
  assign m_2337_io_x1 = m_2191_io_s; // @[MUL.scala 252:21]
  assign m_2337_io_x2 = m_2190_io_cout; // @[MUL.scala 253:22]
  assign m_2337_io_x3 = m_2192_io_out_0; // @[MUL.scala 105:13]
  assign m_2338_io_x1 = m_2193_io_s; // @[MUL.scala 252:21]
  assign m_2338_io_x2 = m_2191_io_cout; // @[MUL.scala 253:22]
  assign m_2338_io_x3 = m_2194_io_out_0; // @[MUL.scala 105:13]
  assign m_2339_io_x1 = m_2195_io_s; // @[MUL.scala 252:21]
  assign m_2339_io_x2 = m_2193_io_cout; // @[MUL.scala 253:22]
  assign m_2339_io_x3 = m_2196_io_out_0; // @[MUL.scala 105:13]
  assign m_2340_io_x1 = m_2197_io_s; // @[MUL.scala 252:21]
  assign m_2340_io_x2 = m_2195_io_cout; // @[MUL.scala 253:22]
  assign m_2340_io_x3 = m_2198_io_out_0; // @[MUL.scala 105:13]
  assign m_2341_io_x1 = m_2199_io_s; // @[MUL.scala 252:21]
  assign m_2341_io_x2 = m_2197_io_cout; // @[MUL.scala 253:22]
  assign m_2341_io_x3 = m_2200_io_out_0; // @[MUL.scala 105:13]
  assign m_2342_io_x1 = m_2201_io_s; // @[MUL.scala 252:21]
  assign m_2342_io_x2 = m_2199_io_cout; // @[MUL.scala 253:22]
  assign m_2342_io_x3 = m_2202_io_out_0; // @[MUL.scala 105:13]
  assign m_2343_io_x1 = m_2203_io_s; // @[MUL.scala 252:21]
  assign m_2343_io_x2 = m_2201_io_cout; // @[MUL.scala 253:22]
  assign m_2343_io_x3 = m_2204_io_out_0; // @[MUL.scala 105:13]
  assign m_2344_io_x1 = m_2205_io_s; // @[MUL.scala 252:21]
  assign m_2344_io_x2 = m_2203_io_cout; // @[MUL.scala 253:22]
  assign m_2344_io_x3 = m_2206_io_out_0; // @[MUL.scala 105:13]
  assign m_2345_io_x1 = m_2207_io_s; // @[MUL.scala 252:21]
  assign m_2345_io_x2 = m_2205_io_cout; // @[MUL.scala 253:22]
  assign m_2345_io_x3 = m_2208_io_out_0; // @[MUL.scala 105:13]
  assign m_2346_io_x1 = m_2209_io_s; // @[MUL.scala 252:21]
  assign m_2346_io_x2 = m_2207_io_cout; // @[MUL.scala 253:22]
  assign m_2346_io_x3 = m_2210_io_out_0; // @[MUL.scala 105:13]
  assign m_2347_io_x1 = m_2211_io_s; // @[MUL.scala 252:21]
  assign m_2347_io_x2 = m_2209_io_cout; // @[MUL.scala 253:22]
  assign m_2347_io_x3 = m_2212_io_out_0; // @[MUL.scala 105:13]
  assign m_2348_io_x1 = m_2213_io_s; // @[MUL.scala 252:21]
  assign m_2348_io_x2 = m_2211_io_cout; // @[MUL.scala 253:22]
  assign m_2348_io_x3 = m_2214_io_out_0; // @[MUL.scala 105:13]
  assign m_2349_io_x1 = m_2215_io_s; // @[MUL.scala 252:21]
  assign m_2349_io_x2 = m_2213_io_cout; // @[MUL.scala 253:22]
  assign m_2349_io_x3 = m_2216_io_out_0; // @[MUL.scala 105:13]
  assign m_2350_io_x1 = m_2217_io_s; // @[MUL.scala 252:21]
  assign m_2350_io_x2 = m_2215_io_cout; // @[MUL.scala 253:22]
  assign m_2350_io_x3 = m_2218_io_out_0; // @[MUL.scala 105:13]
  assign m_2351_io_x1 = m_2219_io_s; // @[MUL.scala 252:21]
  assign m_2351_io_x2 = m_2217_io_cout; // @[MUL.scala 253:22]
  assign m_2351_io_x3 = m_2220_io_out_0; // @[MUL.scala 105:13]
  assign m_2352_io_x1 = m_2221_io_s; // @[MUL.scala 252:21]
  assign m_2352_io_x2 = m_2219_io_cout; // @[MUL.scala 253:22]
  assign m_2352_io_x3 = m_2222_io_out_0; // @[MUL.scala 105:13]
  assign m_2353_io_x1 = m_2223_io_s; // @[MUL.scala 252:21]
  assign m_2353_io_x2 = m_2221_io_cout; // @[MUL.scala 253:22]
  assign m_2353_io_x3 = m_2224_io_out_0; // @[MUL.scala 105:13]
  assign m_2354_io_x1 = m_2225_io_s; // @[MUL.scala 252:21]
  assign m_2354_io_x2 = m_2223_io_cout; // @[MUL.scala 253:22]
  assign m_2354_io_x3 = m_2226_io_out_0; // @[MUL.scala 105:13]
  assign m_2355_io_x1 = m_2227_io_s; // @[MUL.scala 252:21]
  assign m_2355_io_x2 = m_2225_io_cout; // @[MUL.scala 253:22]
  assign m_2355_io_x3 = m_2228_io_out_0; // @[MUL.scala 105:13]
  assign m_2356_io_x1 = m_2229_io_s; // @[MUL.scala 252:21]
  assign m_2356_io_x2 = m_2227_io_cout; // @[MUL.scala 253:22]
  assign m_2356_io_x3 = m_2230_io_out_0; // @[MUL.scala 105:13]
  assign m_2357_io_x1 = m_2231_io_s; // @[MUL.scala 252:21]
  assign m_2357_io_x2 = m_2229_io_cout; // @[MUL.scala 253:22]
  assign m_2357_io_x3 = m_2232_io_out_0; // @[MUL.scala 105:13]
  assign m_2358_io_x1 = m_2233_io_s; // @[MUL.scala 252:21]
  assign m_2358_io_x2 = m_2231_io_cout; // @[MUL.scala 253:22]
  assign m_2358_io_x3 = m_2067_io_cout; // @[MUL.scala 253:22]
  assign m_2359_io_x1 = m_2234_io_s; // @[MUL.scala 252:21]
  assign m_2359_io_x2 = m_2233_io_cout; // @[MUL.scala 253:22]
  assign m_2359_io_x3 = m_2069_io_cout; // @[MUL.scala 253:22]
  assign m_2360_io_x1 = m_2235_io_s; // @[MUL.scala 252:21]
  assign m_2360_io_x2 = m_2234_io_cout; // @[MUL.scala 253:22]
  assign m_2360_io_x3 = m_2071_io_cout; // @[MUL.scala 253:22]
  assign m_2361_io_x1 = m_2236_io_s; // @[MUL.scala 252:21]
  assign m_2361_io_x2 = m_2235_io_cout; // @[MUL.scala 253:22]
  assign m_2361_io_x3 = m_2073_io_cout; // @[MUL.scala 253:22]
  assign m_2362_io_x1 = m_2237_io_s; // @[MUL.scala 252:21]
  assign m_2362_io_x2 = m_2236_io_cout; // @[MUL.scala 253:22]
  assign m_2362_io_x3 = m_2075_io_cout; // @[MUL.scala 253:22]
  assign m_2363_io_x1 = m_2238_io_s; // @[MUL.scala 252:21]
  assign m_2363_io_x2 = m_2237_io_cout; // @[MUL.scala 253:22]
  assign m_2363_io_x3 = m_2077_io_cout; // @[MUL.scala 253:22]
  assign m_2364_io_x1 = m_2239_io_s; // @[MUL.scala 252:21]
  assign m_2364_io_x2 = m_2238_io_cout; // @[MUL.scala 253:22]
  assign m_2364_io_x3 = m_2079_io_cout; // @[MUL.scala 253:22]
  assign m_2365_io_x1 = m_2240_io_s; // @[MUL.scala 252:21]
  assign m_2365_io_x2 = m_2239_io_cout; // @[MUL.scala 253:22]
  assign m_2365_io_x3 = m_2081_io_cout; // @[MUL.scala 253:22]
  assign m_2366_io_x1 = m_2241_io_s; // @[MUL.scala 252:21]
  assign m_2366_io_x2 = m_2240_io_cout; // @[MUL.scala 253:22]
  assign m_2366_io_x3 = m_2083_io_cout; // @[MUL.scala 253:22]
  assign m_2367_io_x1 = m_2242_io_s; // @[MUL.scala 252:21]
  assign m_2367_io_x2 = m_2241_io_cout; // @[MUL.scala 253:22]
  assign m_2367_io_x3 = m_2085_io_cout; // @[MUL.scala 253:22]
  assign m_2368_io_x1 = m_2243_io_s; // @[MUL.scala 252:21]
  assign m_2368_io_x2 = m_2242_io_cout; // @[MUL.scala 253:22]
  assign m_2368_io_x3 = m_2087_io_cout; // @[MUL.scala 253:22]
  assign m_2369_io_x1 = m_2244_io_s; // @[MUL.scala 252:21]
  assign m_2369_io_x2 = m_2243_io_cout; // @[MUL.scala 253:22]
  assign m_2369_io_x3 = m_2089_io_cout; // @[MUL.scala 253:22]
  assign m_2370_io_x1 = m_2245_io_s; // @[MUL.scala 252:21]
  assign m_2370_io_x2 = m_2244_io_cout; // @[MUL.scala 253:22]
  assign m_2370_io_x3 = m_2091_io_cout; // @[MUL.scala 253:22]
  assign m_2371_io_x1 = m_2246_io_s; // @[MUL.scala 252:21]
  assign m_2371_io_x2 = m_2245_io_cout; // @[MUL.scala 253:22]
  assign m_2371_io_x3 = m_2093_io_cout; // @[MUL.scala 253:22]
  assign m_2372_io_x1 = m_2247_io_s; // @[MUL.scala 252:21]
  assign m_2372_io_x2 = m_2246_io_cout; // @[MUL.scala 253:22]
  assign m_2372_io_x3 = m_2095_io_out_1; // @[MUL.scala 105:13]
  assign m_2373_io_x1 = m_2248_io_s; // @[MUL.scala 252:21]
  assign m_2373_io_x2 = m_2247_io_cout; // @[MUL.scala 253:22]
  assign m_2373_io_x3 = m_2097_io_out_1; // @[MUL.scala 105:13]
  assign m_2374_io_x1 = m_2249_io_s; // @[MUL.scala 252:21]
  assign m_2374_io_x2 = m_2248_io_cout; // @[MUL.scala 253:22]
  assign m_2374_io_x3 = m_2099_io_out_1; // @[MUL.scala 105:13]
  assign m_2375_io_x1 = m_2250_io_s; // @[MUL.scala 252:21]
  assign m_2375_io_x2 = m_2249_io_cout; // @[MUL.scala 253:22]
  assign m_2375_io_x3 = m_2101_io_out_1; // @[MUL.scala 105:13]
  assign m_2376_io_x1 = m_2251_io_s; // @[MUL.scala 252:21]
  assign m_2376_io_x2 = m_2250_io_cout; // @[MUL.scala 253:22]
  assign m_2376_io_x3 = m_2103_io_out_1; // @[MUL.scala 105:13]
  assign m_2377_io_in_0 = m_2252_io_s; // @[MUL.scala 252:21]
  assign m_2377_io_in_1 = m_2251_io_cout; // @[MUL.scala 253:22]
  assign m_2378_io_in_0 = m_2253_io_s; // @[MUL.scala 252:21]
  assign m_2378_io_in_1 = m_2252_io_cout; // @[MUL.scala 253:22]
  assign m_2379_io_in_0 = m_2254_io_s; // @[MUL.scala 252:21]
  assign m_2379_io_in_1 = m_2253_io_cout; // @[MUL.scala 253:22]
  assign m_2380_io_in_0 = m_2255_io_s; // @[MUL.scala 252:21]
  assign m_2380_io_in_1 = m_2254_io_cout; // @[MUL.scala 253:22]
  assign m_2381_io_in_0 = m_2256_io_s; // @[MUL.scala 252:21]
  assign m_2381_io_in_1 = m_2255_io_cout; // @[MUL.scala 253:22]
  assign m_2382_io_in_0 = m_2257_io_s; // @[MUL.scala 252:21]
  assign m_2382_io_in_1 = m_2256_io_cout; // @[MUL.scala 253:22]
  assign m_2383_io_in_0 = m_2258_io_s; // @[MUL.scala 252:21]
  assign m_2383_io_in_1 = m_2257_io_cout; // @[MUL.scala 253:22]
  assign m_2384_io_in_0 = m_2259_io_s; // @[MUL.scala 252:21]
  assign m_2384_io_in_1 = m_2258_io_cout; // @[MUL.scala 253:22]
  assign m_2385_io_in_0 = m_2260_io_s; // @[MUL.scala 252:21]
  assign m_2385_io_in_1 = m_2259_io_cout; // @[MUL.scala 253:22]
  assign m_2386_io_in_0 = m_2261_io_s; // @[MUL.scala 252:21]
  assign m_2386_io_in_1 = m_2260_io_cout; // @[MUL.scala 253:22]
  assign m_2387_io_in_0 = m_2262_io_s; // @[MUL.scala 252:21]
  assign m_2387_io_in_1 = m_2261_io_cout; // @[MUL.scala 253:22]
  assign m_2388_io_in_0 = m_2263_io_out_0; // @[MUL.scala 125:16]
  assign m_2388_io_in_1 = m_2262_io_cout; // @[MUL.scala 253:22]
  assign m_2389_io_in_0 = m_2264_io_out_0; // @[MUL.scala 125:16]
  assign m_2389_io_in_1 = m_2263_io_out_1; // @[MUL.scala 126:16]
  assign m_2390_io_in_0 = m_2265_io_out_0; // @[MUL.scala 125:16]
  assign m_2390_io_in_1 = m_2264_io_out_1; // @[MUL.scala 126:16]
  assign m_2391_io_in_0 = m_2266_io_out_0; // @[MUL.scala 125:16]
  assign m_2391_io_in_1 = m_2265_io_out_1; // @[MUL.scala 126:16]
  assign m_2392_io_in_0 = m_2267_io_out_0; // @[MUL.scala 125:16]
  assign m_2392_io_in_1 = m_2266_io_out_1; // @[MUL.scala 126:16]
  assign m_2393_io_in_0 = m_2268_io_out_0; // @[MUL.scala 125:16]
  assign m_2393_io_in_1 = m_2267_io_out_1; // @[MUL.scala 126:16]
  assign m_2394_io_in_0 = m_2269_io_out_0; // @[MUL.scala 125:16]
  assign m_2394_io_in_1 = m_2268_io_out_1; // @[MUL.scala 126:16]
  assign m_2395_io_in_0 = m_2270_io_out_0; // @[MUL.scala 125:16]
  assign m_2395_io_in_1 = m_2269_io_out_1; // @[MUL.scala 126:16]
  assign m_2396_io_in_0 = m_2271_io_out_0; // @[MUL.scala 125:16]
  assign m_2396_io_in_1 = m_2270_io_out_1; // @[MUL.scala 126:16]
  assign m_2397_io_in_0 = m_2272_io_out_0; // @[MUL.scala 125:16]
  assign m_2397_io_in_1 = m_2271_io_out_1; // @[MUL.scala 126:16]
  assign m_2398_io_in_0 = m_2273_io_out_0; // @[MUL.scala 125:16]
  assign m_2398_io_in_1 = m_2272_io_out_1; // @[MUL.scala 126:16]
  assign m_2399_io_in_0 = m_2274_io_out_0; // @[MUL.scala 125:16]
  assign m_2399_io_in_1 = m_2273_io_out_1; // @[MUL.scala 126:16]
  assign m_2400_io_in_0 = m_2275_io_out_0; // @[MUL.scala 125:16]
  assign m_2400_io_in_1 = m_2274_io_out_1; // @[MUL.scala 126:16]
  assign m_2401_io_in_0 = m_2276_io_out_0; // @[MUL.scala 125:16]
  assign m_2401_io_in_1 = m_2275_io_out_1; // @[MUL.scala 126:16]
  assign m_2402_io_in_0 = m_2277_io_out_0; // @[MUL.scala 125:16]
  assign m_2402_io_in_1 = m_2276_io_out_1; // @[MUL.scala 126:16]
  assign m_2403_io_in_0 = m_2278_io_out_0; // @[MUL.scala 125:16]
  assign m_2403_io_in_1 = m_2277_io_out_1; // @[MUL.scala 126:16]
  assign m_2404_io_in_0 = m_2279_io_out_0; // @[MUL.scala 125:16]
  assign m_2404_io_in_1 = m_2278_io_out_1; // @[MUL.scala 126:16]
  assign m_2405_io_in_0 = m_2280_io_out_0; // @[MUL.scala 125:16]
  assign m_2405_io_in_1 = m_2279_io_out_1; // @[MUL.scala 126:16]
  assign m_2406_io_in_0 = m_2281_io_out_0; // @[MUL.scala 125:16]
  assign m_2406_io_in_1 = m_2280_io_out_1; // @[MUL.scala 126:16]
  assign m_2407_io_in_0 = m_2282_io_out_0; // @[MUL.scala 125:16]
  assign m_2407_io_in_1 = m_2281_io_out_1; // @[MUL.scala 126:16]
  assign m_2408_io_in_0 = m_2283_io_out_0; // @[MUL.scala 125:16]
  assign m_2408_io_in_1 = m_2282_io_out_1; // @[MUL.scala 126:16]
  assign m_2409_io_in_0 = m_2284_io_out_0; // @[MUL.scala 125:16]
  assign m_2409_io_in_1 = m_2283_io_out_1; // @[MUL.scala 126:16]
  assign m_2410_io_in_0 = m_2285_io_out_0; // @[MUL.scala 125:16]
  assign m_2410_io_in_1 = m_2284_io_out_1; // @[MUL.scala 126:16]
  assign m_2411_io_in_0 = m_2287_io_out_0; // @[MUL.scala 125:16]
  assign m_2411_io_in_1 = m_2286_io_out_1; // @[MUL.scala 126:16]
  assign m_2412_io_in_0 = m_2288_io_out_0; // @[MUL.scala 125:16]
  assign m_2412_io_in_1 = m_2287_io_out_1; // @[MUL.scala 126:16]
  assign m_2413_io_in_0 = m_2289_io_out_0; // @[MUL.scala 125:16]
  assign m_2413_io_in_1 = m_2288_io_out_1; // @[MUL.scala 126:16]
  assign m_2414_io_in_0 = m_2290_io_out_0; // @[MUL.scala 125:16]
  assign m_2414_io_in_1 = m_2289_io_out_1; // @[MUL.scala 126:16]
  assign m_2415_io_in_0 = m_2291_io_out_0; // @[MUL.scala 125:16]
  assign m_2415_io_in_1 = m_2290_io_out_1; // @[MUL.scala 126:16]
  assign m_2416_io_in_0 = m_2292_io_out_0; // @[MUL.scala 125:16]
  assign m_2416_io_in_1 = m_2291_io_out_1; // @[MUL.scala 126:16]
  assign m_2417_io_in_0 = m_2293_io_out_0; // @[MUL.scala 125:16]
  assign m_2417_io_in_1 = m_2292_io_out_1; // @[MUL.scala 126:16]
  assign m_2418_io_in_0 = m_2294_io_out_0; // @[MUL.scala 125:16]
  assign m_2418_io_in_1 = m_2293_io_out_1; // @[MUL.scala 126:16]
  assign m_2419_io_in_0 = m_2295_io_out_0; // @[MUL.scala 125:16]
  assign m_2419_io_in_1 = m_2294_io_out_1; // @[MUL.scala 126:16]
  assign m_2420_io_in_0 = m_2296_io_out_0; // @[MUL.scala 125:16]
  assign m_2420_io_in_1 = m_2295_io_out_1; // @[MUL.scala 126:16]
  assign m_2421_io_in_0 = m_2297_io_out_0; // @[MUL.scala 125:16]
  assign m_2421_io_in_1 = m_2296_io_out_1; // @[MUL.scala 126:16]
  assign m_2422_io_in_0 = m_2298_io_out_0; // @[MUL.scala 125:16]
  assign m_2422_io_in_1 = m_2297_io_out_1; // @[MUL.scala 126:16]
  assign m_2423_io_in_0 = m_2299_io_out_0; // @[MUL.scala 125:16]
  assign m_2423_io_in_1 = m_2298_io_out_1; // @[MUL.scala 126:16]
  assign m_2424_io_in_0 = m_2300_io_out_0; // @[MUL.scala 125:16]
  assign m_2424_io_in_1 = m_2299_io_out_1; // @[MUL.scala 126:16]
  assign m_2425_io_in_0 = m_2301_io_out_0; // @[MUL.scala 125:16]
  assign m_2425_io_in_1 = m_2300_io_out_1; // @[MUL.scala 126:16]
  assign m_2426_io_in_0 = m_2302_io_out_0; // @[MUL.scala 125:16]
  assign m_2426_io_in_1 = m_2301_io_out_1; // @[MUL.scala 126:16]
  assign m_2427_io_in_0 = m_2303_io_out_0; // @[MUL.scala 125:16]
  assign m_2427_io_in_1 = m_2302_io_out_1; // @[MUL.scala 126:16]
  assign m_2428_io_in_0 = m_2304_io_out_0; // @[MUL.scala 125:16]
  assign m_2428_io_in_1 = m_2303_io_out_1; // @[MUL.scala 126:16]
  assign m_2429_io_in_0 = m_2305_io_out_0; // @[MUL.scala 125:16]
  assign m_2429_io_in_1 = m_2304_io_out_1; // @[MUL.scala 126:16]
  assign m_2430_io_in_0 = m_2306_io_out_0; // @[MUL.scala 125:16]
  assign m_2430_io_in_1 = m_2305_io_out_1; // @[MUL.scala 126:16]
  assign m_2431_io_in_0 = m_2307_io_out_0; // @[MUL.scala 125:16]
  assign m_2431_io_in_1 = m_2306_io_out_1; // @[MUL.scala 126:16]
  assign m_2432_io_in_0 = m_2308_io_out_0; // @[MUL.scala 125:16]
  assign m_2432_io_in_1 = m_2307_io_out_1; // @[MUL.scala 126:16]
  assign m_2433_io_in_0 = m_2309_io_out_0; // @[MUL.scala 125:16]
  assign m_2433_io_in_1 = m_2308_io_out_1; // @[MUL.scala 126:16]
  assign m_2434_io_in_0 = m_2310_io_out_0; // @[MUL.scala 125:16]
  assign m_2434_io_in_1 = m_2309_io_out_1; // @[MUL.scala 126:16]
  assign m_2435_io_in_0 = m_2311_io_out_0; // @[MUL.scala 125:16]
  assign m_2435_io_in_1 = m_2310_io_out_1; // @[MUL.scala 126:16]
  assign m_2436_io_in_0 = m_2312_io_out_0; // @[MUL.scala 125:16]
  assign m_2436_io_in_1 = m_2311_io_out_1; // @[MUL.scala 126:16]
  assign m_2437_io_in_0 = m_2313_io_out_0; // @[MUL.scala 125:16]
  assign m_2437_io_in_1 = m_2312_io_out_1; // @[MUL.scala 126:16]
  assign m_2438_io_in_0 = m_2314_io_out_0; // @[MUL.scala 125:16]
  assign m_2438_io_in_1 = m_2313_io_out_1; // @[MUL.scala 126:16]
  assign m_2439_io_in_0 = m_2315_io_out_0; // @[MUL.scala 125:16]
  assign m_2439_io_in_1 = m_2314_io_out_1; // @[MUL.scala 126:16]
  assign m_2440_io_in_0 = m_2316_io_out_0; // @[MUL.scala 125:16]
  assign m_2440_io_in_1 = m_2315_io_out_1; // @[MUL.scala 126:16]
  assign m_2441_io_in_0 = m_2317_io_out_0; // @[MUL.scala 125:16]
  assign m_2441_io_in_1 = m_2316_io_out_1; // @[MUL.scala 126:16]
  assign m_2442_io_in_0 = m_2318_io_out_0; // @[MUL.scala 125:16]
  assign m_2442_io_in_1 = m_2317_io_out_1; // @[MUL.scala 126:16]
  assign m_2443_io_in_0 = m_2319_io_s; // @[MUL.scala 252:21]
  assign m_2443_io_in_1 = m_2318_io_out_1; // @[MUL.scala 126:16]
  assign m_2444_io_in_0 = m_2320_io_s; // @[MUL.scala 252:21]
  assign m_2444_io_in_1 = m_2319_io_cout; // @[MUL.scala 253:22]
  assign m_2445_io_in_0 = m_2321_io_s; // @[MUL.scala 252:21]
  assign m_2445_io_in_1 = m_2320_io_cout; // @[MUL.scala 253:22]
  assign m_2446_io_in_0 = m_2322_io_s; // @[MUL.scala 252:21]
  assign m_2446_io_in_1 = m_2321_io_cout; // @[MUL.scala 253:22]
  assign m_2447_io_in_0 = m_2323_io_s; // @[MUL.scala 252:21]
  assign m_2447_io_in_1 = m_2322_io_cout; // @[MUL.scala 253:22]
  assign m_2448_io_in_0 = m_2324_io_s; // @[MUL.scala 252:21]
  assign m_2448_io_in_1 = m_2323_io_cout; // @[MUL.scala 253:22]
  assign m_2449_io_in_0 = m_2325_io_s; // @[MUL.scala 252:21]
  assign m_2449_io_in_1 = m_2324_io_cout; // @[MUL.scala 253:22]
  assign m_2450_io_in_0 = m_2326_io_s; // @[MUL.scala 252:21]
  assign m_2450_io_in_1 = m_2325_io_cout; // @[MUL.scala 253:22]
  assign m_2451_io_in_0 = m_2327_io_s; // @[MUL.scala 252:21]
  assign m_2451_io_in_1 = m_2326_io_cout; // @[MUL.scala 253:22]
  assign m_2452_io_in_0 = m_2328_io_s; // @[MUL.scala 252:21]
  assign m_2452_io_in_1 = m_2327_io_cout; // @[MUL.scala 253:22]
  assign m_2453_io_in_0 = m_2329_io_s; // @[MUL.scala 252:21]
  assign m_2453_io_in_1 = m_2328_io_cout; // @[MUL.scala 253:22]
  assign m_2454_io_in_0 = m_2330_io_s; // @[MUL.scala 252:21]
  assign m_2454_io_in_1 = m_2329_io_cout; // @[MUL.scala 253:22]
  assign m_2455_io_in_0 = m_2331_io_s; // @[MUL.scala 252:21]
  assign m_2455_io_in_1 = m_2330_io_cout; // @[MUL.scala 253:22]
  assign m_2456_io_in_0 = m_2332_io_s; // @[MUL.scala 252:21]
  assign m_2456_io_in_1 = m_2331_io_cout; // @[MUL.scala 253:22]
  assign m_2457_io_in_0 = m_2333_io_s; // @[MUL.scala 252:21]
  assign m_2457_io_in_1 = m_2332_io_cout; // @[MUL.scala 253:22]
  assign m_2458_io_in_0 = m_2334_io_s; // @[MUL.scala 252:21]
  assign m_2458_io_in_1 = m_2333_io_cout; // @[MUL.scala 253:22]
  assign m_2459_io_in_0 = m_2335_io_s; // @[MUL.scala 252:21]
  assign m_2459_io_in_1 = m_2334_io_cout; // @[MUL.scala 253:22]
  assign m_2460_io_in_0 = m_2336_io_s; // @[MUL.scala 252:21]
  assign m_2460_io_in_1 = m_2335_io_cout; // @[MUL.scala 253:22]
  assign m_2461_io_in_0 = m_2337_io_s; // @[MUL.scala 252:21]
  assign m_2461_io_in_1 = m_2336_io_cout; // @[MUL.scala 253:22]
  assign m_2462_io_x1 = m_2338_io_s; // @[MUL.scala 252:21]
  assign m_2462_io_x2 = m_2337_io_cout; // @[MUL.scala 253:22]
  assign m_2462_io_x3 = m_2192_io_out_1; // @[MUL.scala 105:13]
  assign m_2463_io_x1 = m_2339_io_s; // @[MUL.scala 252:21]
  assign m_2463_io_x2 = m_2338_io_cout; // @[MUL.scala 253:22]
  assign m_2463_io_x3 = m_2194_io_out_1; // @[MUL.scala 105:13]
  assign m_2464_io_x1 = m_2340_io_s; // @[MUL.scala 252:21]
  assign m_2464_io_x2 = m_2339_io_cout; // @[MUL.scala 253:22]
  assign m_2464_io_x3 = m_2196_io_out_1; // @[MUL.scala 105:13]
  assign m_2465_io_x1 = m_2341_io_s; // @[MUL.scala 252:21]
  assign m_2465_io_x2 = m_2340_io_cout; // @[MUL.scala 253:22]
  assign m_2465_io_x3 = m_2198_io_out_1; // @[MUL.scala 105:13]
  assign m_2466_io_x1 = m_2342_io_s; // @[MUL.scala 252:21]
  assign m_2466_io_x2 = m_2341_io_cout; // @[MUL.scala 253:22]
  assign m_2466_io_x3 = m_2200_io_out_1; // @[MUL.scala 105:13]
  assign m_2467_io_x1 = m_2343_io_s; // @[MUL.scala 252:21]
  assign m_2467_io_x2 = m_2342_io_cout; // @[MUL.scala 253:22]
  assign m_2467_io_x3 = m_2202_io_out_1; // @[MUL.scala 105:13]
  assign m_2468_io_x1 = m_2344_io_s; // @[MUL.scala 252:21]
  assign m_2468_io_x2 = m_2343_io_cout; // @[MUL.scala 253:22]
  assign m_2468_io_x3 = m_2204_io_out_1; // @[MUL.scala 105:13]
  assign m_2469_io_x1 = m_2345_io_s; // @[MUL.scala 252:21]
  assign m_2469_io_x2 = m_2344_io_cout; // @[MUL.scala 253:22]
  assign m_2469_io_x3 = m_2206_io_out_1; // @[MUL.scala 105:13]
  assign m_2470_io_x1 = m_2346_io_s; // @[MUL.scala 252:21]
  assign m_2470_io_x2 = m_2345_io_cout; // @[MUL.scala 253:22]
  assign m_2470_io_x3 = m_2208_io_out_1; // @[MUL.scala 105:13]
  assign m_2471_io_x1 = m_2347_io_s; // @[MUL.scala 252:21]
  assign m_2471_io_x2 = m_2346_io_cout; // @[MUL.scala 253:22]
  assign m_2471_io_x3 = m_2210_io_out_1; // @[MUL.scala 105:13]
  assign m_2472_io_x1 = m_2348_io_s; // @[MUL.scala 252:21]
  assign m_2472_io_x2 = m_2347_io_cout; // @[MUL.scala 253:22]
  assign m_2472_io_x3 = m_2212_io_out_1; // @[MUL.scala 105:13]
  assign m_2473_io_x1 = m_2349_io_s; // @[MUL.scala 252:21]
  assign m_2473_io_x2 = m_2348_io_cout; // @[MUL.scala 253:22]
  assign m_2473_io_x3 = m_2214_io_out_1; // @[MUL.scala 105:13]
  assign m_2474_io_x1 = m_2350_io_s; // @[MUL.scala 252:21]
  assign m_2474_io_x2 = m_2349_io_cout; // @[MUL.scala 253:22]
  assign m_2474_io_x3 = m_2216_io_out_1; // @[MUL.scala 105:13]
  assign m_2475_io_x1 = m_2351_io_s; // @[MUL.scala 252:21]
  assign m_2475_io_x2 = m_2350_io_cout; // @[MUL.scala 253:22]
  assign m_2475_io_x3 = m_2218_io_out_1; // @[MUL.scala 105:13]
  assign m_2476_io_x1 = m_2352_io_s; // @[MUL.scala 252:21]
  assign m_2476_io_x2 = m_2351_io_cout; // @[MUL.scala 253:22]
  assign m_2476_io_x3 = m_2220_io_out_1; // @[MUL.scala 105:13]
  assign m_2477_io_x1 = m_2353_io_s; // @[MUL.scala 252:21]
  assign m_2477_io_x2 = m_2352_io_cout; // @[MUL.scala 253:22]
  assign m_2477_io_x3 = m_2222_io_out_1; // @[MUL.scala 105:13]
  assign m_2478_io_x1 = m_2354_io_s; // @[MUL.scala 252:21]
  assign m_2478_io_x2 = m_2353_io_cout; // @[MUL.scala 253:22]
  assign m_2478_io_x3 = m_2224_io_out_1; // @[MUL.scala 105:13]
  assign m_2479_io_x1 = m_2355_io_s; // @[MUL.scala 252:21]
  assign m_2479_io_x2 = m_2354_io_cout; // @[MUL.scala 253:22]
  assign m_2479_io_x3 = m_2226_io_out_1; // @[MUL.scala 105:13]
  assign m_2480_io_x1 = m_2356_io_s; // @[MUL.scala 252:21]
  assign m_2480_io_x2 = m_2355_io_cout; // @[MUL.scala 253:22]
  assign m_2480_io_x3 = m_2228_io_out_1; // @[MUL.scala 105:13]
  assign m_2481_io_x1 = m_2357_io_s; // @[MUL.scala 252:21]
  assign m_2481_io_x2 = m_2356_io_cout; // @[MUL.scala 253:22]
  assign m_2481_io_x3 = m_2230_io_out_1; // @[MUL.scala 105:13]
  assign m_2482_io_x1 = m_2358_io_s; // @[MUL.scala 252:21]
  assign m_2482_io_x2 = m_2357_io_cout; // @[MUL.scala 253:22]
  assign m_2482_io_x3 = m_2232_io_out_1; // @[MUL.scala 105:13]
  assign m_2483_io_in_0 = m_2359_io_s; // @[MUL.scala 252:21]
  assign m_2483_io_in_1 = m_2358_io_cout; // @[MUL.scala 253:22]
  assign m_2484_io_in_0 = m_2360_io_s; // @[MUL.scala 252:21]
  assign m_2484_io_in_1 = m_2359_io_cout; // @[MUL.scala 253:22]
  assign m_2485_io_in_0 = m_2361_io_s; // @[MUL.scala 252:21]
  assign m_2485_io_in_1 = m_2360_io_cout; // @[MUL.scala 253:22]
  assign m_2486_io_in_0 = m_2362_io_s; // @[MUL.scala 252:21]
  assign m_2486_io_in_1 = m_2361_io_cout; // @[MUL.scala 253:22]
  assign m_2487_io_in_0 = m_2363_io_s; // @[MUL.scala 252:21]
  assign m_2487_io_in_1 = m_2362_io_cout; // @[MUL.scala 253:22]
  assign m_2488_io_in_0 = m_2364_io_s; // @[MUL.scala 252:21]
  assign m_2488_io_in_1 = m_2363_io_cout; // @[MUL.scala 253:22]
  assign m_2489_io_in_0 = m_2365_io_s; // @[MUL.scala 252:21]
  assign m_2489_io_in_1 = m_2364_io_cout; // @[MUL.scala 253:22]
  assign m_2490_io_in_0 = m_2366_io_s; // @[MUL.scala 252:21]
  assign m_2490_io_in_1 = m_2365_io_cout; // @[MUL.scala 253:22]
  assign m_2491_io_in_0 = m_2367_io_s; // @[MUL.scala 252:21]
  assign m_2491_io_in_1 = m_2366_io_cout; // @[MUL.scala 253:22]
  assign m_2492_io_in_0 = m_2368_io_s; // @[MUL.scala 252:21]
  assign m_2492_io_in_1 = m_2367_io_cout; // @[MUL.scala 253:22]
  assign m_2493_io_in_0 = m_2369_io_s; // @[MUL.scala 252:21]
  assign m_2493_io_in_1 = m_2368_io_cout; // @[MUL.scala 253:22]
  assign m_2494_io_in_0 = m_2370_io_s; // @[MUL.scala 252:21]
  assign m_2494_io_in_1 = m_2369_io_cout; // @[MUL.scala 253:22]
  assign m_2495_io_in_0 = m_2371_io_s; // @[MUL.scala 252:21]
  assign m_2495_io_in_1 = m_2370_io_cout; // @[MUL.scala 253:22]
  assign m_2496_io_in_0 = m_2372_io_s; // @[MUL.scala 252:21]
  assign m_2496_io_in_1 = m_2371_io_cout; // @[MUL.scala 253:22]
  assign m_2497_io_in_0 = m_2373_io_s; // @[MUL.scala 252:21]
  assign m_2497_io_in_1 = m_2372_io_cout; // @[MUL.scala 253:22]
  assign m_2498_io_in_0 = m_2374_io_s; // @[MUL.scala 252:21]
  assign m_2498_io_in_1 = m_2373_io_cout; // @[MUL.scala 253:22]
  assign m_2499_io_in_0 = m_2375_io_s; // @[MUL.scala 252:21]
  assign m_2499_io_in_1 = m_2374_io_cout; // @[MUL.scala 253:22]
  assign m_2500_io_in_0 = m_2376_io_s; // @[MUL.scala 252:21]
  assign m_2500_io_in_1 = m_2375_io_cout; // @[MUL.scala 253:22]
  assign m_2501_io_in_0 = m_2377_io_out_0; // @[MUL.scala 125:16]
  assign m_2501_io_in_1 = m_2376_io_cout; // @[MUL.scala 253:22]
  assign m_2502_io_in_0 = m_2378_io_out_0; // @[MUL.scala 125:16]
  assign m_2502_io_in_1 = m_2377_io_out_1; // @[MUL.scala 126:16]
  assign m_2503_io_in_0 = m_2379_io_out_0; // @[MUL.scala 125:16]
  assign m_2503_io_in_1 = m_2378_io_out_1; // @[MUL.scala 126:16]
  assign m_2504_io_in_0 = m_2380_io_out_0; // @[MUL.scala 125:16]
  assign m_2504_io_in_1 = m_2379_io_out_1; // @[MUL.scala 126:16]
  assign m_2505_io_in_0 = m_2381_io_out_0; // @[MUL.scala 125:16]
  assign m_2505_io_in_1 = m_2380_io_out_1; // @[MUL.scala 126:16]
  assign m_2506_io_in_0 = m_2382_io_out_0; // @[MUL.scala 125:16]
  assign m_2506_io_in_1 = m_2381_io_out_1; // @[MUL.scala 126:16]
  assign m_2507_io_in_0 = m_2383_io_out_0; // @[MUL.scala 125:16]
  assign m_2507_io_in_1 = m_2382_io_out_1; // @[MUL.scala 126:16]
  assign m_2508_io_in_0 = m_2384_io_out_0; // @[MUL.scala 125:16]
  assign m_2508_io_in_1 = m_2383_io_out_1; // @[MUL.scala 126:16]
  assign m_2509_io_in_0 = m_2385_io_out_0; // @[MUL.scala 125:16]
  assign m_2509_io_in_1 = m_2384_io_out_1; // @[MUL.scala 126:16]
  assign m_2510_io_in_0 = m_2386_io_out_0; // @[MUL.scala 125:16]
  assign m_2510_io_in_1 = m_2385_io_out_1; // @[MUL.scala 126:16]
  assign m_2511_io_in_0 = m_2387_io_out_0; // @[MUL.scala 125:16]
  assign m_2511_io_in_1 = m_2386_io_out_1; // @[MUL.scala 126:16]
  assign m_2512_io_in_0 = m_2388_io_out_0; // @[MUL.scala 125:16]
  assign m_2512_io_in_1 = m_2387_io_out_1; // @[MUL.scala 126:16]
  assign m_2513_io_in_0 = m_2389_io_out_0; // @[MUL.scala 125:16]
  assign m_2513_io_in_1 = m_2388_io_out_1; // @[MUL.scala 126:16]
  assign m_2514_io_in_0 = m_2390_io_out_0; // @[MUL.scala 125:16]
  assign m_2514_io_in_1 = m_2389_io_out_1; // @[MUL.scala 126:16]
  assign m_2515_io_in_0 = m_2391_io_out_0; // @[MUL.scala 125:16]
  assign m_2515_io_in_1 = m_2390_io_out_1; // @[MUL.scala 126:16]
  assign m_2516_io_in_0 = m_2392_io_out_0; // @[MUL.scala 125:16]
  assign m_2516_io_in_1 = m_2391_io_out_1; // @[MUL.scala 126:16]
  assign m_2517_io_in_0 = m_2393_io_out_0; // @[MUL.scala 125:16]
  assign m_2517_io_in_1 = m_2392_io_out_1; // @[MUL.scala 126:16]
  assign m_2518_io_in_0 = m_2394_io_out_0; // @[MUL.scala 125:16]
  assign m_2518_io_in_1 = m_2393_io_out_1; // @[MUL.scala 126:16]
  assign m_2519_io_in_0 = m_2395_io_out_0; // @[MUL.scala 125:16]
  assign m_2519_io_in_1 = m_2394_io_out_1; // @[MUL.scala 126:16]
  assign m_2520_io_in_0 = m_2396_io_out_0; // @[MUL.scala 125:16]
  assign m_2520_io_in_1 = m_2395_io_out_1; // @[MUL.scala 126:16]
  assign m_2521_io_in_0 = m_2397_io_out_0; // @[MUL.scala 125:16]
  assign m_2521_io_in_1 = m_2396_io_out_1; // @[MUL.scala 126:16]
  assign m_2522_io_in_0 = m_2398_io_out_0; // @[MUL.scala 125:16]
  assign m_2522_io_in_1 = m_2397_io_out_1; // @[MUL.scala 126:16]
  assign m_2523_io_in_0 = m_2399_io_out_0; // @[MUL.scala 125:16]
  assign m_2523_io_in_1 = m_2398_io_out_1; // @[MUL.scala 126:16]
  assign m_2524_io_in_0 = m_2400_io_out_0; // @[MUL.scala 125:16]
  assign m_2524_io_in_1 = m_2399_io_out_1; // @[MUL.scala 126:16]
  assign m_2525_io_in_0 = m_2401_io_out_0; // @[MUL.scala 125:16]
  assign m_2525_io_in_1 = m_2400_io_out_1; // @[MUL.scala 126:16]
  assign m_2526_io_in_0 = m_2402_io_out_0; // @[MUL.scala 125:16]
  assign m_2526_io_in_1 = m_2401_io_out_1; // @[MUL.scala 126:16]
  assign m_2527_io_in_0 = m_2403_io_out_0; // @[MUL.scala 125:16]
  assign m_2527_io_in_1 = m_2402_io_out_1; // @[MUL.scala 126:16]
  assign m_2528_io_in_0 = m_2404_io_out_0; // @[MUL.scala 125:16]
  assign m_2528_io_in_1 = m_2403_io_out_1; // @[MUL.scala 126:16]
  assign m_2529_io_in_0 = m_2405_io_out_0; // @[MUL.scala 125:16]
  assign m_2529_io_in_1 = m_2404_io_out_1; // @[MUL.scala 126:16]
  assign m_2530_io_in_0 = m_2406_io_out_0; // @[MUL.scala 125:16]
  assign m_2530_io_in_1 = m_2405_io_out_1; // @[MUL.scala 126:16]
  assign m_2531_io_in_0 = m_2407_io_out_0; // @[MUL.scala 125:16]
  assign m_2531_io_in_1 = m_2406_io_out_1; // @[MUL.scala 126:16]
  assign m_2532_io_in_0 = m_2408_io_out_0; // @[MUL.scala 125:16]
  assign m_2532_io_in_1 = m_2407_io_out_1; // @[MUL.scala 126:16]
  assign m_2533_io_in_0 = m_2409_io_out_0; // @[MUL.scala 125:16]
  assign m_2533_io_in_1 = m_2408_io_out_1; // @[MUL.scala 126:16]
  assign m_2534_io_in_0 = m_2410_io_out_0; // @[MUL.scala 125:16]
  assign m_2534_io_in_1 = m_2409_io_out_1; // @[MUL.scala 126:16]
  always @(posedge clock) begin
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r <= m_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1 <= m_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2 <= m_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_3 <= m_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_4 <= m_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_5 <= m_1_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_6 <= m_1_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_7 <= m_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_8 <= m_1_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_9 <= m_1_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_10 <= m_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_11 <= m_1_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_12 <= m_2_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_13 <= m_2_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_14 <= m_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_15 <= m_1_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_16 <= m_2_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_17 <= m_2_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_18 <= m_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_19 <= m_1_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_20 <= m_2_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_21 <= m_3_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_22 <= m_3_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_23 <= m_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_24 <= m_1_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_25 <= m_2_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_26 <= m_3_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_27 <= m_3_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_28 <= m_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_29 <= m_1_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_30 <= m_2_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_31 <= m_3_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_32 <= m_4_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_33 <= m_4_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_34 <= m_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_35 <= m_1_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_36 <= m_2_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_37 <= m_3_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_38 <= m_4_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_39 <= m_4_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_40 <= m_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_41 <= m_1_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_42 <= m_2_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_43 <= m_3_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_44 <= m_4_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_45 <= m_5_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_46 <= m_5_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_47 <= m_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_48 <= m_1_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_49 <= m_2_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_50 <= m_3_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_51 <= m_4_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_52 <= m_5_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_53 <= m_5_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_54 <= m_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_55 <= m_1_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_56 <= m_2_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_57 <= m_3_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_58 <= m_4_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_59 <= m_5_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_60 <= m_6_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_61 <= m_6_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_62 <= m_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_63 <= m_1_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_64 <= m_2_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_65 <= m_3_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_66 <= m_4_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_67 <= m_5_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_68 <= m_6_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_69 <= m_6_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_70 <= m_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_71 <= m_1_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_72 <= m_2_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_73 <= m_3_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_74 <= m_4_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_75 <= m_5_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_76 <= m_6_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_77 <= m_7_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_78 <= m_7_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_79 <= m_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_80 <= m_1_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_81 <= m_2_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_82 <= m_3_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_83 <= m_4_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_84 <= m_5_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_85 <= m_6_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_86 <= m_7_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_87 <= m_7_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_88 <= m_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_89 <= m_1_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_90 <= m_2_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_91 <= m_3_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_92 <= m_4_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_93 <= m_5_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_94 <= m_6_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_95 <= m_7_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_96 <= m_8_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_97 <= m_8_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_98 <= m_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_99 <= m_1_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_100 <= m_2_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_101 <= m_3_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_102 <= m_4_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_103 <= m_5_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_104 <= m_6_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_105 <= m_7_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_106 <= m_8_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_107 <= m_8_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_108 <= m_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_109 <= m_1_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_110 <= m_2_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_111 <= m_3_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_112 <= m_4_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_113 <= m_5_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_114 <= m_6_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_115 <= m_7_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_116 <= m_8_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_117 <= m_9_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_118 <= m_9_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_119 <= m_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_120 <= m_1_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_121 <= m_2_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_122 <= m_3_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_123 <= m_4_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_124 <= m_5_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_125 <= m_6_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_126 <= m_7_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_127 <= m_8_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_128 <= m_9_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_129 <= m_9_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_130 <= m_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_131 <= m_1_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_132 <= m_2_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_133 <= m_3_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_134 <= m_4_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_135 <= m_5_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_136 <= m_6_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_137 <= m_7_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_138 <= m_8_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_139 <= m_9_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_140 <= m_10_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_141 <= m_10_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_142 <= m_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_143 <= m_1_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_144 <= m_2_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_145 <= m_3_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_146 <= m_4_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_147 <= m_5_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_148 <= m_6_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_149 <= m_7_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_150 <= m_8_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_151 <= m_9_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_152 <= m_10_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_153 <= m_10_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_154 <= m_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_155 <= m_1_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_156 <= m_2_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_157 <= m_3_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_158 <= m_4_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_159 <= m_5_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_160 <= m_6_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_161 <= m_7_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_162 <= m_8_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_163 <= m_9_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_164 <= m_10_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_165 <= m_11_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_166 <= m_11_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_167 <= m_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_168 <= m_1_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_169 <= m_2_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_170 <= m_3_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_171 <= m_4_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_172 <= m_5_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_173 <= m_6_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_174 <= m_7_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_175 <= m_8_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_176 <= m_9_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_177 <= m_10_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_178 <= m_11_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_179 <= m_11_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_180 <= m_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_181 <= m_1_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_182 <= m_2_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_183 <= m_3_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_184 <= m_4_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_185 <= m_5_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_186 <= m_6_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_187 <= m_7_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_188 <= m_8_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_189 <= m_9_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_190 <= m_10_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_191 <= m_11_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_192 <= m_12_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_193 <= m_12_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_194 <= m_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_195 <= m_1_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_196 <= m_2_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_197 <= m_3_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_198 <= m_4_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_199 <= m_5_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_200 <= m_6_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_201 <= m_7_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_202 <= m_8_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_203 <= m_9_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_204 <= m_10_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_205 <= m_11_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_206 <= m_12_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_207 <= m_12_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_208 <= m_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_209 <= m_1_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_210 <= m_2_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_211 <= m_3_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_212 <= m_4_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_213 <= m_5_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_214 <= m_6_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_215 <= m_7_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_216 <= m_8_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_217 <= m_9_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_218 <= m_10_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_219 <= m_11_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_220 <= m_12_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_221 <= m_13_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_222 <= m_13_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_223 <= m_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_224 <= m_1_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_225 <= m_2_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_226 <= m_3_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_227 <= m_4_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_228 <= m_5_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_229 <= m_6_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_230 <= m_7_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_231 <= m_8_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_232 <= m_9_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_233 <= m_10_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_234 <= m_11_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_235 <= m_12_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_236 <= m_13_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_237 <= m_13_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_238 <= m_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_239 <= m_1_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_240 <= m_2_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_241 <= m_3_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_242 <= m_4_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_243 <= m_5_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_244 <= m_6_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_245 <= m_7_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_246 <= m_8_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_247 <= m_9_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_248 <= m_10_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_249 <= m_11_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_250 <= m_12_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_251 <= m_13_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_252 <= m_14_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_253 <= m_14_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_254 <= m_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_255 <= m_1_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_256 <= m_2_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_257 <= m_3_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_258 <= m_4_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_259 <= m_5_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_260 <= m_6_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_261 <= m_7_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_262 <= m_8_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_263 <= m_9_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_264 <= m_10_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_265 <= m_11_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_266 <= m_12_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_267 <= m_13_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_268 <= m_14_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_269 <= m_14_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_270 <= m_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_271 <= m_1_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_272 <= m_2_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_273 <= m_3_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_274 <= m_4_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_275 <= m_5_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_276 <= m_6_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_277 <= m_7_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_278 <= m_8_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_279 <= m_9_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_280 <= m_10_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_281 <= m_11_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_282 <= m_12_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_283 <= m_13_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_284 <= m_14_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_285 <= m_15_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_286 <= m_15_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_287 <= m_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_288 <= m_1_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_289 <= m_2_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_290 <= m_3_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_291 <= m_4_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_292 <= m_5_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_293 <= m_6_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_294 <= m_7_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_295 <= m_8_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_296 <= m_9_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_297 <= m_10_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_298 <= m_11_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_299 <= m_12_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_300 <= m_13_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_301 <= m_14_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_302 <= m_15_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_303 <= m_15_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_304 <= m_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_305 <= m_1_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_306 <= m_2_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_307 <= m_3_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_308 <= m_4_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_309 <= m_5_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_310 <= m_6_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_311 <= m_7_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_312 <= m_8_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_313 <= m_9_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_314 <= m_10_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_315 <= m_11_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_316 <= m_12_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_317 <= m_13_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_318 <= m_14_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_319 <= m_15_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_320 <= m_16_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_321 <= m_16_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_322 <= m_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_323 <= m_1_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_324 <= m_2_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_325 <= m_3_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_326 <= m_4_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_327 <= m_5_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_328 <= m_6_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_329 <= m_7_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_330 <= m_8_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_331 <= m_9_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_332 <= m_10_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_333 <= m_11_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_334 <= m_12_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_335 <= m_13_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_336 <= m_14_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_337 <= m_15_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_338 <= m_16_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_339 <= m_16_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_340 <= m_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_341 <= m_1_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_342 <= m_2_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_343 <= m_3_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_344 <= m_4_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_345 <= m_5_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_346 <= m_6_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_347 <= m_7_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_348 <= m_8_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_349 <= m_9_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_350 <= m_10_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_351 <= m_11_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_352 <= m_12_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_353 <= m_13_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_354 <= m_14_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_355 <= m_15_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_356 <= m_16_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_357 <= m_17_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_358 <= m_17_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_359 <= m_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_360 <= m_1_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_361 <= m_2_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_362 <= m_3_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_363 <= m_4_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_364 <= m_5_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_365 <= m_6_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_366 <= m_7_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_367 <= m_8_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_368 <= m_9_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_369 <= m_10_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_370 <= m_11_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_371 <= m_12_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_372 <= m_13_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_373 <= m_14_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_374 <= m_15_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_375 <= m_16_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_376 <= m_17_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_377 <= m_17_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_378 <= m_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_379 <= m_1_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_380 <= m_2_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_381 <= m_3_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_382 <= m_4_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_383 <= m_5_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_384 <= m_6_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_385 <= m_7_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_386 <= m_8_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_387 <= m_9_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_388 <= m_10_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_389 <= m_11_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_390 <= m_12_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_391 <= m_13_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_392 <= m_14_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_393 <= m_15_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_394 <= m_16_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_395 <= m_17_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_396 <= m_18_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_397 <= m_18_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_398 <= m_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_399 <= m_1_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_400 <= m_2_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_401 <= m_3_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_402 <= m_4_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_403 <= m_5_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_404 <= m_6_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_405 <= m_7_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_406 <= m_8_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_407 <= m_9_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_408 <= m_10_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_409 <= m_11_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_410 <= m_12_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_411 <= m_13_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_412 <= m_14_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_413 <= m_15_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_414 <= m_16_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_415 <= m_17_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_416 <= m_18_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_417 <= m_18_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_418 <= m_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_419 <= m_1_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_420 <= m_2_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_421 <= m_3_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_422 <= m_4_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_423 <= m_5_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_424 <= m_6_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_425 <= m_7_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_426 <= m_8_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_427 <= m_9_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_428 <= m_10_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_429 <= m_11_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_430 <= m_12_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_431 <= m_13_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_432 <= m_14_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_433 <= m_15_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_434 <= m_16_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_435 <= m_17_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_436 <= m_18_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_437 <= m_19_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_438 <= m_19_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_439 <= m_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_440 <= m_1_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_441 <= m_2_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_442 <= m_3_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_443 <= m_4_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_444 <= m_5_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_445 <= m_6_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_446 <= m_7_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_447 <= m_8_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_448 <= m_9_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_449 <= m_10_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_450 <= m_11_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_451 <= m_12_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_452 <= m_13_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_453 <= m_14_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_454 <= m_15_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_455 <= m_16_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_456 <= m_17_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_457 <= m_18_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_458 <= m_19_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_459 <= m_19_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_460 <= m_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_461 <= m_1_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_462 <= m_2_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_463 <= m_3_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_464 <= m_4_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_465 <= m_5_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_466 <= m_6_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_467 <= m_7_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_468 <= m_8_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_469 <= m_9_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_470 <= m_10_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_471 <= m_11_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_472 <= m_12_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_473 <= m_13_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_474 <= m_14_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_475 <= m_15_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_476 <= m_16_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_477 <= m_17_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_478 <= m_18_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_479 <= m_19_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_480 <= m_20_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_481 <= m_20_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_482 <= m_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_483 <= m_1_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_484 <= m_2_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_485 <= m_3_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_486 <= m_4_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_487 <= m_5_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_488 <= m_6_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_489 <= m_7_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_490 <= m_8_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_491 <= m_9_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_492 <= m_10_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_493 <= m_11_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_494 <= m_12_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_495 <= m_13_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_496 <= m_14_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_497 <= m_15_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_498 <= m_16_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_499 <= m_17_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_500 <= m_18_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_501 <= m_19_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_502 <= m_20_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_503 <= m_20_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_504 <= m_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_505 <= m_1_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_506 <= m_2_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_507 <= m_3_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_508 <= m_4_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_509 <= m_5_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_510 <= m_6_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_511 <= m_7_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_512 <= m_8_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_513 <= m_9_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_514 <= m_10_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_515 <= m_11_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_516 <= m_12_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_517 <= m_13_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_518 <= m_14_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_519 <= m_15_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_520 <= m_16_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_521 <= m_17_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_522 <= m_18_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_523 <= m_19_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_524 <= m_20_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_525 <= m_21_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_526 <= m_21_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_527 <= m_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_528 <= m_1_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_529 <= m_2_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_530 <= m_3_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_531 <= m_4_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_532 <= m_5_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_533 <= m_6_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_534 <= m_7_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_535 <= m_8_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_536 <= m_9_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_537 <= m_10_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_538 <= m_11_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_539 <= m_12_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_540 <= m_13_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_541 <= m_14_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_542 <= m_15_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_543 <= m_16_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_544 <= m_17_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_545 <= m_18_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_546 <= m_19_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_547 <= m_20_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_548 <= m_21_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_549 <= m_21_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_550 <= m_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_551 <= m_1_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_552 <= m_2_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_553 <= m_3_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_554 <= m_4_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_555 <= m_5_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_556 <= m_6_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_557 <= m_7_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_558 <= m_8_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_559 <= m_9_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_560 <= m_10_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_561 <= m_11_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_562 <= m_12_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_563 <= m_13_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_564 <= m_14_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_565 <= m_15_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_566 <= m_16_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_567 <= m_17_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_568 <= m_18_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_569 <= m_19_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_570 <= m_20_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_571 <= m_21_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_572 <= m_22_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_573 <= m_22_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_574 <= m_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_575 <= m_1_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_576 <= m_2_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_577 <= m_3_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_578 <= m_4_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_579 <= m_5_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_580 <= m_6_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_581 <= m_7_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_582 <= m_8_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_583 <= m_9_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_584 <= m_10_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_585 <= m_11_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_586 <= m_12_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_587 <= m_13_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_588 <= m_14_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_589 <= m_15_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_590 <= m_16_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_591 <= m_17_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_592 <= m_18_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_593 <= m_19_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_594 <= m_20_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_595 <= m_21_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_596 <= m_22_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_597 <= m_22_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_598 <= m_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_599 <= m_1_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_600 <= m_2_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_601 <= m_3_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_602 <= m_4_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_603 <= m_5_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_604 <= m_6_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_605 <= m_7_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_606 <= m_8_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_607 <= m_9_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_608 <= m_10_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_609 <= m_11_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_610 <= m_12_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_611 <= m_13_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_612 <= m_14_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_613 <= m_15_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_614 <= m_16_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_615 <= m_17_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_616 <= m_18_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_617 <= m_19_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_618 <= m_20_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_619 <= m_21_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_620 <= m_22_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_621 <= m_23_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_622 <= m_23_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_623 <= m_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_624 <= m_1_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_625 <= m_2_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_626 <= m_3_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_627 <= m_4_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_628 <= m_5_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_629 <= m_6_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_630 <= m_7_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_631 <= m_8_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_632 <= m_9_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_633 <= m_10_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_634 <= m_11_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_635 <= m_12_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_636 <= m_13_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_637 <= m_14_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_638 <= m_15_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_639 <= m_16_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_640 <= m_17_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_641 <= m_18_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_642 <= m_19_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_643 <= m_20_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_644 <= m_21_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_645 <= m_22_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_646 <= m_23_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_647 <= m_23_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_648 <= m_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_649 <= m_1_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_650 <= m_2_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_651 <= m_3_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_652 <= m_4_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_653 <= m_5_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_654 <= m_6_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_655 <= m_7_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_656 <= m_8_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_657 <= m_9_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_658 <= m_10_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_659 <= m_11_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_660 <= m_12_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_661 <= m_13_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_662 <= m_14_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_663 <= m_15_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_664 <= m_16_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_665 <= m_17_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_666 <= m_18_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_667 <= m_19_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_668 <= m_20_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_669 <= m_21_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_670 <= m_22_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_671 <= m_23_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_672 <= m_24_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_673 <= m_24_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_674 <= m_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_675 <= m_1_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_676 <= m_2_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_677 <= m_3_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_678 <= m_4_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_679 <= m_5_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_680 <= m_6_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_681 <= m_7_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_682 <= m_8_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_683 <= m_9_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_684 <= m_10_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_685 <= m_11_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_686 <= m_12_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_687 <= m_13_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_688 <= m_14_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_689 <= m_15_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_690 <= m_16_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_691 <= m_17_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_692 <= m_18_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_693 <= m_19_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_694 <= m_20_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_695 <= m_21_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_696 <= m_22_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_697 <= m_23_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_698 <= m_24_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_699 <= m_24_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_700 <= m_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_701 <= m_1_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_702 <= m_2_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_703 <= m_3_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_704 <= m_4_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_705 <= m_5_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_706 <= m_6_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_707 <= m_7_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_708 <= m_8_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_709 <= m_9_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_710 <= m_10_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_711 <= m_11_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_712 <= m_12_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_713 <= m_13_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_714 <= m_14_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_715 <= m_15_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_716 <= m_16_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_717 <= m_17_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_718 <= m_18_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_719 <= m_19_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_720 <= m_20_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_721 <= m_21_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_722 <= m_22_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_723 <= m_23_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_724 <= m_24_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_725 <= m_25_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_726 <= m_25_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_727 <= m_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_728 <= m_1_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_729 <= m_2_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_730 <= m_3_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_731 <= m_4_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_732 <= m_5_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_733 <= m_6_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_734 <= m_7_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_735 <= m_8_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_736 <= m_9_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_737 <= m_10_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_738 <= m_11_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_739 <= m_12_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_740 <= m_13_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_741 <= m_14_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_742 <= m_15_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_743 <= m_16_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_744 <= m_17_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_745 <= m_18_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_746 <= m_19_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_747 <= m_20_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_748 <= m_21_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_749 <= m_22_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_750 <= m_23_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_751 <= m_24_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_752 <= m_25_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_753 <= m_25_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_754 <= m_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_755 <= m_1_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_756 <= m_2_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_757 <= m_3_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_758 <= m_4_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_759 <= m_5_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_760 <= m_6_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_761 <= m_7_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_762 <= m_8_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_763 <= m_9_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_764 <= m_10_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_765 <= m_11_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_766 <= m_12_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_767 <= m_13_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_768 <= m_14_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_769 <= m_15_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_770 <= m_16_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_771 <= m_17_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_772 <= m_18_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_773 <= m_19_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_774 <= m_20_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_775 <= m_21_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_776 <= m_22_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_777 <= m_23_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_778 <= m_24_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_779 <= m_25_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_780 <= m_26_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_781 <= m_26_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_782 <= m_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_783 <= m_1_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_784 <= m_2_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_785 <= m_3_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_786 <= m_4_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_787 <= m_5_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_788 <= m_6_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_789 <= m_7_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_790 <= m_8_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_791 <= m_9_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_792 <= m_10_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_793 <= m_11_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_794 <= m_12_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_795 <= m_13_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_796 <= m_14_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_797 <= m_15_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_798 <= m_16_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_799 <= m_17_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_800 <= m_18_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_801 <= m_19_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_802 <= m_20_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_803 <= m_21_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_804 <= m_22_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_805 <= m_23_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_806 <= m_24_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_807 <= m_25_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_808 <= m_26_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_809 <= m_26_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_810 <= m_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_811 <= m_1_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_812 <= m_2_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_813 <= m_3_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_814 <= m_4_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_815 <= m_5_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_816 <= m_6_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_817 <= m_7_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_818 <= m_8_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_819 <= m_9_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_820 <= m_10_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_821 <= m_11_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_822 <= m_12_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_823 <= m_13_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_824 <= m_14_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_825 <= m_15_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_826 <= m_16_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_827 <= m_17_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_828 <= m_18_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_829 <= m_19_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_830 <= m_20_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_831 <= m_21_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_832 <= m_22_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_833 <= m_23_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_834 <= m_24_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_835 <= m_25_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_836 <= m_26_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_837 <= m_27_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_838 <= m_27_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_839 <= m_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_840 <= m_1_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_841 <= m_2_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_842 <= m_3_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_843 <= m_4_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_844 <= m_5_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_845 <= m_6_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_846 <= m_7_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_847 <= m_8_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_848 <= m_9_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_849 <= m_10_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_850 <= m_11_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_851 <= m_12_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_852 <= m_13_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_853 <= m_14_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_854 <= m_15_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_855 <= m_16_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_856 <= m_17_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_857 <= m_18_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_858 <= m_19_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_859 <= m_20_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_860 <= m_21_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_861 <= m_22_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_862 <= m_23_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_863 <= m_24_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_864 <= m_25_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_865 <= m_26_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_866 <= m_27_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_867 <= m_27_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_868 <= m_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_869 <= m_1_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_870 <= m_2_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_871 <= m_3_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_872 <= m_4_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_873 <= m_5_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_874 <= m_6_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_875 <= m_7_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_876 <= m_8_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_877 <= m_9_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_878 <= m_10_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_879 <= m_11_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_880 <= m_12_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_881 <= m_13_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_882 <= m_14_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_883 <= m_15_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_884 <= m_16_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_885 <= m_17_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_886 <= m_18_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_887 <= m_19_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_888 <= m_20_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_889 <= m_21_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_890 <= m_22_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_891 <= m_23_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_892 <= m_24_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_893 <= m_25_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_894 <= m_26_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_895 <= m_27_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_896 <= m_28_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_897 <= m_28_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_898 <= m_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_899 <= m_1_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_900 <= m_2_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_901 <= m_3_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_902 <= m_4_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_903 <= m_5_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_904 <= m_6_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_905 <= m_7_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_906 <= m_8_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_907 <= m_9_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_908 <= m_10_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_909 <= m_11_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_910 <= m_12_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_911 <= m_13_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_912 <= m_14_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_913 <= m_15_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_914 <= m_16_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_915 <= m_17_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_916 <= m_18_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_917 <= m_19_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_918 <= m_20_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_919 <= m_21_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_920 <= m_22_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_921 <= m_23_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_922 <= m_24_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_923 <= m_25_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_924 <= m_26_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_925 <= m_27_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_926 <= m_28_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_927 <= m_28_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_928 <= m_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_929 <= m_1_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_930 <= m_2_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_931 <= m_3_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_932 <= m_4_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_933 <= m_5_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_934 <= m_6_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_935 <= m_7_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_936 <= m_8_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_937 <= m_9_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_938 <= m_10_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_939 <= m_11_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_940 <= m_12_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_941 <= m_13_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_942 <= m_14_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_943 <= m_15_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_944 <= m_16_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_945 <= m_17_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_946 <= m_18_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_947 <= m_19_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_948 <= m_20_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_949 <= m_21_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_950 <= m_22_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_951 <= m_23_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_952 <= m_24_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_953 <= m_25_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_954 <= m_26_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_955 <= m_27_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_956 <= m_28_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_957 <= m_29_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_958 <= m_29_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_959 <= m_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_960 <= m_1_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_961 <= m_2_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_962 <= m_3_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_963 <= m_4_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_964 <= m_5_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_965 <= m_6_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_966 <= m_7_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_967 <= m_8_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_968 <= m_9_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_969 <= m_10_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_970 <= m_11_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_971 <= m_12_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_972 <= m_13_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_973 <= m_14_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_974 <= m_15_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_975 <= m_16_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_976 <= m_17_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_977 <= m_18_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_978 <= m_19_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_979 <= m_20_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_980 <= m_21_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_981 <= m_22_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_982 <= m_23_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_983 <= m_24_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_984 <= m_25_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_985 <= m_26_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_986 <= m_27_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_987 <= m_28_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_988 <= m_29_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_989 <= m_29_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_990 <= m_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_991 <= m_1_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_992 <= m_2_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_993 <= m_3_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_994 <= m_4_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_995 <= m_5_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_996 <= m_6_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_997 <= m_7_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_998 <= m_8_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_999 <= m_9_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1000 <= m_10_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1001 <= m_11_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1002 <= m_12_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1003 <= m_13_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1004 <= m_14_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1005 <= m_15_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1006 <= m_16_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1007 <= m_17_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1008 <= m_18_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1009 <= m_19_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1010 <= m_20_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1011 <= m_21_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1012 <= m_22_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1013 <= m_23_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1014 <= m_24_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1015 <= m_25_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1016 <= m_26_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1017 <= m_27_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1018 <= m_28_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1019 <= m_29_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1020 <= m_30_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1021 <= m_30_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1022 <= m_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1023 <= m_1_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1024 <= m_2_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1025 <= m_3_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1026 <= m_4_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1027 <= m_5_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1028 <= m_6_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1029 <= m_7_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1030 <= m_8_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1031 <= m_9_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1032 <= m_10_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1033 <= m_11_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1034 <= m_12_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1035 <= m_13_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1036 <= m_14_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1037 <= m_15_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1038 <= m_16_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1039 <= m_17_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1040 <= m_18_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1041 <= m_19_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1042 <= m_20_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1043 <= m_21_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1044 <= m_22_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1045 <= m_23_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1046 <= m_24_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1047 <= m_25_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1048 <= m_26_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1049 <= m_27_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1050 <= m_28_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1051 <= m_29_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1052 <= m_30_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1053 <= m_30_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1054 <= m_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1055 <= m_1_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1056 <= m_2_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1057 <= m_3_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1058 <= m_4_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1059 <= m_5_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1060 <= m_6_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1061 <= m_7_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1062 <= m_8_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1063 <= m_9_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1064 <= m_10_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1065 <= m_11_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1066 <= m_12_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1067 <= m_13_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1068 <= m_14_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1069 <= m_15_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1070 <= m_16_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1071 <= m_17_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1072 <= m_18_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1073 <= m_19_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1074 <= m_20_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1075 <= m_21_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1076 <= m_22_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1077 <= m_23_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1078 <= m_24_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1079 <= m_25_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1080 <= m_26_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1081 <= m_27_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1082 <= m_28_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1083 <= m_29_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1084 <= m_30_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1085 <= m_31_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1086 <= m_31_io_carry[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1087 <= m_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1088 <= m_1_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1089 <= m_2_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1090 <= m_3_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1091 <= m_4_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1092 <= m_5_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1093 <= m_6_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1094 <= m_7_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1095 <= m_8_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1096 <= m_9_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1097 <= m_10_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1098 <= m_11_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1099 <= m_12_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1100 <= m_13_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1101 <= m_14_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1102 <= m_15_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1103 <= m_16_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1104 <= m_17_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1105 <= m_18_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1106 <= m_19_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1107 <= m_20_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1108 <= m_21_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1109 <= m_22_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1110 <= m_23_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1111 <= m_24_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1112 <= m_25_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1113 <= m_26_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1114 <= m_27_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1115 <= m_28_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1116 <= m_29_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1117 <= m_30_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1118 <= m_31_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1119 <= m_31_io_carry[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1120 <= m_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1121 <= m_1_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1122 <= m_2_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1123 <= m_3_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1124 <= m_4_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1125 <= m_5_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1126 <= m_6_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1127 <= m_7_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1128 <= m_8_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1129 <= m_9_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1130 <= m_10_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1131 <= m_11_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1132 <= m_12_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1133 <= m_13_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1134 <= m_14_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1135 <= m_15_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1136 <= m_16_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1137 <= m_17_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1138 <= m_18_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1139 <= m_19_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1140 <= m_20_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1141 <= m_21_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1142 <= m_22_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1143 <= m_23_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1144 <= m_24_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1145 <= m_25_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1146 <= m_26_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1147 <= m_27_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1148 <= m_28_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1149 <= m_29_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1150 <= m_30_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1151 <= m_31_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1152 <= m_32_io_p[0]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1153 <= m_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1154 <= m_1_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1155 <= m_2_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1156 <= m_3_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1157 <= m_4_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1158 <= m_5_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1159 <= m_6_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1160 <= m_7_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1161 <= m_8_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1162 <= m_9_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1163 <= m_10_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1164 <= m_11_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1165 <= m_12_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1166 <= m_13_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1167 <= m_14_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1168 <= m_15_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1169 <= m_16_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1170 <= m_17_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1171 <= m_18_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1172 <= m_19_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1173 <= m_20_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1174 <= m_21_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1175 <= m_22_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1176 <= m_23_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1177 <= m_24_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1178 <= m_25_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1179 <= m_26_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1180 <= m_27_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1181 <= m_28_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1182 <= m_29_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1183 <= m_30_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1184 <= m_31_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1185 <= m_32_io_p[1]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1186 <= m_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1187 <= m_1_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1188 <= m_2_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1189 <= m_3_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1190 <= m_4_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1191 <= m_5_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1192 <= m_6_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1193 <= m_7_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1194 <= m_8_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1195 <= m_9_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1196 <= m_10_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1197 <= m_11_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1198 <= m_12_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1199 <= m_13_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1200 <= m_14_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1201 <= m_15_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1202 <= m_16_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1203 <= m_17_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1204 <= m_18_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1205 <= m_19_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1206 <= m_20_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1207 <= m_21_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1208 <= m_22_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1209 <= m_23_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1210 <= m_24_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1211 <= m_25_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1212 <= m_26_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1213 <= m_27_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1214 <= m_28_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1215 <= m_29_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1216 <= m_30_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1217 <= m_31_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1218 <= m_32_io_p[2]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1219 <= m_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1220 <= m_1_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1221 <= m_2_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1222 <= m_3_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1223 <= m_4_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1224 <= m_5_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1225 <= m_6_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1226 <= m_7_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1227 <= m_8_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1228 <= m_9_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1229 <= m_10_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1230 <= m_11_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1231 <= m_12_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1232 <= m_13_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1233 <= m_14_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1234 <= m_15_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1235 <= m_16_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1236 <= m_17_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1237 <= m_18_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1238 <= m_19_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1239 <= m_20_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1240 <= m_21_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1241 <= m_22_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1242 <= m_23_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1243 <= m_24_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1244 <= m_25_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1245 <= m_26_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1246 <= m_27_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1247 <= m_28_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1248 <= m_29_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1249 <= m_30_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1250 <= m_31_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1251 <= m_32_io_p[3]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1252 <= _T_88; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1253 <= _T_157; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1254 <= m_2_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1255 <= m_3_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1256 <= m_4_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1257 <= m_5_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1258 <= m_6_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1259 <= m_7_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1260 <= m_8_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1261 <= m_9_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1262 <= m_10_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1263 <= m_11_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1264 <= m_12_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1265 <= m_13_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1266 <= m_14_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1267 <= m_15_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1268 <= m_16_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1269 <= m_17_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1270 <= m_18_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1271 <= m_19_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1272 <= m_20_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1273 <= m_21_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1274 <= m_22_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1275 <= m_23_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1276 <= m_24_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1277 <= m_25_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1278 <= m_26_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1279 <= m_27_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1280 <= m_28_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1281 <= m_29_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1282 <= m_30_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1283 <= m_31_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1284 <= m_32_io_p[4]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1286 <= m_2_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1287 <= m_3_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1288 <= m_4_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1289 <= m_5_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1290 <= m_6_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1291 <= m_7_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1292 <= m_8_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1293 <= m_9_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1294 <= m_10_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1295 <= m_11_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1296 <= m_12_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1297 <= m_13_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1298 <= m_14_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1299 <= m_15_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1300 <= m_16_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1301 <= m_17_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1302 <= m_18_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1303 <= m_19_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1304 <= m_20_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1305 <= m_21_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1306 <= m_22_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1307 <= m_23_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1308 <= m_24_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1309 <= m_25_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1310 <= m_26_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1311 <= m_27_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1312 <= m_28_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1313 <= m_29_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1314 <= m_30_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1315 <= m_31_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1316 <= m_32_io_p[5]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1317 <= _T_228; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1318 <= m_3_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1319 <= m_4_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1320 <= m_5_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1321 <= m_6_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1322 <= m_7_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1323 <= m_8_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1324 <= m_9_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1325 <= m_10_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1326 <= m_11_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1327 <= m_12_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1328 <= m_13_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1329 <= m_14_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1330 <= m_15_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1331 <= m_16_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1332 <= m_17_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1333 <= m_18_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1334 <= m_19_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1335 <= m_20_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1336 <= m_21_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1337 <= m_22_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1338 <= m_23_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1339 <= m_24_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1340 <= m_25_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1341 <= m_26_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1342 <= m_27_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1343 <= m_28_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1344 <= m_29_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1345 <= m_30_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1346 <= m_31_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1347 <= m_32_io_p[6]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1349 <= m_3_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1350 <= m_4_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1351 <= m_5_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1352 <= m_6_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1353 <= m_7_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1354 <= m_8_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1355 <= m_9_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1356 <= m_10_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1357 <= m_11_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1358 <= m_12_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1359 <= m_13_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1360 <= m_14_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1361 <= m_15_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1362 <= m_16_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1363 <= m_17_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1364 <= m_18_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1365 <= m_19_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1366 <= m_20_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1367 <= m_21_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1368 <= m_22_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1369 <= m_23_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1370 <= m_24_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1371 <= m_25_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1372 <= m_26_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1373 <= m_27_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1374 <= m_28_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1375 <= m_29_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1376 <= m_30_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1377 <= m_31_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1378 <= m_32_io_p[7]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1379 <= _T_299; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1380 <= m_4_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1381 <= m_5_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1382 <= m_6_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1383 <= m_7_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1384 <= m_8_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1385 <= m_9_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1386 <= m_10_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1387 <= m_11_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1388 <= m_12_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1389 <= m_13_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1390 <= m_14_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1391 <= m_15_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1392 <= m_16_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1393 <= m_17_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1394 <= m_18_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1395 <= m_19_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1396 <= m_20_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1397 <= m_21_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1398 <= m_22_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1399 <= m_23_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1400 <= m_24_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1401 <= m_25_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1402 <= m_26_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1403 <= m_27_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1404 <= m_28_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1405 <= m_29_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1406 <= m_30_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1407 <= m_31_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1408 <= m_32_io_p[8]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1410 <= m_4_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1411 <= m_5_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1412 <= m_6_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1413 <= m_7_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1414 <= m_8_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1415 <= m_9_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1416 <= m_10_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1417 <= m_11_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1418 <= m_12_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1419 <= m_13_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1420 <= m_14_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1421 <= m_15_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1422 <= m_16_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1423 <= m_17_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1424 <= m_18_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1425 <= m_19_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1426 <= m_20_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1427 <= m_21_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1428 <= m_22_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1429 <= m_23_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1430 <= m_24_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1431 <= m_25_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1432 <= m_26_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1433 <= m_27_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1434 <= m_28_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1435 <= m_29_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1436 <= m_30_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1437 <= m_31_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1438 <= m_32_io_p[9]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1439 <= _T_370; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1440 <= m_5_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1441 <= m_6_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1442 <= m_7_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1443 <= m_8_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1444 <= m_9_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1445 <= m_10_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1446 <= m_11_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1447 <= m_12_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1448 <= m_13_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1449 <= m_14_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1450 <= m_15_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1451 <= m_16_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1452 <= m_17_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1453 <= m_18_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1454 <= m_19_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1455 <= m_20_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1456 <= m_21_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1457 <= m_22_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1458 <= m_23_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1459 <= m_24_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1460 <= m_25_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1461 <= m_26_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1462 <= m_27_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1463 <= m_28_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1464 <= m_29_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1465 <= m_30_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1466 <= m_31_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1467 <= m_32_io_p[10]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1469 <= m_5_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1470 <= m_6_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1471 <= m_7_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1472 <= m_8_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1473 <= m_9_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1474 <= m_10_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1475 <= m_11_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1476 <= m_12_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1477 <= m_13_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1478 <= m_14_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1479 <= m_15_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1480 <= m_16_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1481 <= m_17_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1482 <= m_18_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1483 <= m_19_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1484 <= m_20_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1485 <= m_21_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1486 <= m_22_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1487 <= m_23_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1488 <= m_24_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1489 <= m_25_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1490 <= m_26_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1491 <= m_27_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1492 <= m_28_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1493 <= m_29_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1494 <= m_30_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1495 <= m_31_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1496 <= m_32_io_p[11]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1497 <= _T_441; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1498 <= m_6_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1499 <= m_7_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1500 <= m_8_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1501 <= m_9_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1502 <= m_10_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1503 <= m_11_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1504 <= m_12_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1505 <= m_13_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1506 <= m_14_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1507 <= m_15_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1508 <= m_16_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1509 <= m_17_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1510 <= m_18_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1511 <= m_19_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1512 <= m_20_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1513 <= m_21_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1514 <= m_22_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1515 <= m_23_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1516 <= m_24_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1517 <= m_25_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1518 <= m_26_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1519 <= m_27_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1520 <= m_28_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1521 <= m_29_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1522 <= m_30_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1523 <= m_31_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1524 <= m_32_io_p[12]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1526 <= m_6_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1527 <= m_7_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1528 <= m_8_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1529 <= m_9_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1530 <= m_10_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1531 <= m_11_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1532 <= m_12_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1533 <= m_13_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1534 <= m_14_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1535 <= m_15_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1536 <= m_16_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1537 <= m_17_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1538 <= m_18_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1539 <= m_19_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1540 <= m_20_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1541 <= m_21_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1542 <= m_22_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1543 <= m_23_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1544 <= m_24_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1545 <= m_25_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1546 <= m_26_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1547 <= m_27_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1548 <= m_28_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1549 <= m_29_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1550 <= m_30_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1551 <= m_31_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1552 <= m_32_io_p[13]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1553 <= _T_512; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1554 <= m_7_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1555 <= m_8_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1556 <= m_9_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1557 <= m_10_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1558 <= m_11_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1559 <= m_12_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1560 <= m_13_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1561 <= m_14_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1562 <= m_15_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1563 <= m_16_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1564 <= m_17_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1565 <= m_18_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1566 <= m_19_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1567 <= m_20_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1568 <= m_21_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1569 <= m_22_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1570 <= m_23_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1571 <= m_24_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1572 <= m_25_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1573 <= m_26_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1574 <= m_27_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1575 <= m_28_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1576 <= m_29_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1577 <= m_30_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1578 <= m_31_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1579 <= m_32_io_p[14]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1581 <= m_7_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1582 <= m_8_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1583 <= m_9_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1584 <= m_10_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1585 <= m_11_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1586 <= m_12_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1587 <= m_13_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1588 <= m_14_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1589 <= m_15_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1590 <= m_16_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1591 <= m_17_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1592 <= m_18_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1593 <= m_19_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1594 <= m_20_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1595 <= m_21_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1596 <= m_22_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1597 <= m_23_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1598 <= m_24_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1599 <= m_25_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1600 <= m_26_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1601 <= m_27_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1602 <= m_28_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1603 <= m_29_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1604 <= m_30_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1605 <= m_31_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1606 <= m_32_io_p[15]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1607 <= _T_583; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1608 <= m_8_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1609 <= m_9_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1610 <= m_10_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1611 <= m_11_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1612 <= m_12_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1613 <= m_13_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1614 <= m_14_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1615 <= m_15_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1616 <= m_16_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1617 <= m_17_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1618 <= m_18_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1619 <= m_19_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1620 <= m_20_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1621 <= m_21_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1622 <= m_22_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1623 <= m_23_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1624 <= m_24_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1625 <= m_25_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1626 <= m_26_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1627 <= m_27_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1628 <= m_28_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1629 <= m_29_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1630 <= m_30_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1631 <= m_31_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1632 <= m_32_io_p[16]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1634 <= m_8_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1635 <= m_9_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1636 <= m_10_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1637 <= m_11_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1638 <= m_12_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1639 <= m_13_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1640 <= m_14_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1641 <= m_15_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1642 <= m_16_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1643 <= m_17_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1644 <= m_18_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1645 <= m_19_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1646 <= m_20_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1647 <= m_21_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1648 <= m_22_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1649 <= m_23_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1650 <= m_24_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1651 <= m_25_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1652 <= m_26_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1653 <= m_27_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1654 <= m_28_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1655 <= m_29_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1656 <= m_30_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1657 <= m_31_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1658 <= m_32_io_p[17]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1659 <= _T_654; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1660 <= m_9_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1661 <= m_10_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1662 <= m_11_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1663 <= m_12_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1664 <= m_13_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1665 <= m_14_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1666 <= m_15_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1667 <= m_16_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1668 <= m_17_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1669 <= m_18_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1670 <= m_19_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1671 <= m_20_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1672 <= m_21_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1673 <= m_22_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1674 <= m_23_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1675 <= m_24_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1676 <= m_25_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1677 <= m_26_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1678 <= m_27_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1679 <= m_28_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1680 <= m_29_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1681 <= m_30_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1682 <= m_31_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1683 <= m_32_io_p[18]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1685 <= m_9_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1686 <= m_10_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1687 <= m_11_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1688 <= m_12_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1689 <= m_13_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1690 <= m_14_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1691 <= m_15_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1692 <= m_16_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1693 <= m_17_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1694 <= m_18_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1695 <= m_19_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1696 <= m_20_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1697 <= m_21_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1698 <= m_22_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1699 <= m_23_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1700 <= m_24_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1701 <= m_25_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1702 <= m_26_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1703 <= m_27_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1704 <= m_28_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1705 <= m_29_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1706 <= m_30_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1707 <= m_31_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1708 <= m_32_io_p[19]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1709 <= _T_725; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1710 <= m_10_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1711 <= m_11_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1712 <= m_12_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1713 <= m_13_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1714 <= m_14_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1715 <= m_15_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1716 <= m_16_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1717 <= m_17_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1718 <= m_18_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1719 <= m_19_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1720 <= m_20_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1721 <= m_21_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1722 <= m_22_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1723 <= m_23_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1724 <= m_24_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1725 <= m_25_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1726 <= m_26_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1727 <= m_27_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1728 <= m_28_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1729 <= m_29_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1730 <= m_30_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1731 <= m_31_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1732 <= m_32_io_p[20]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1734 <= m_10_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1735 <= m_11_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1736 <= m_12_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1737 <= m_13_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1738 <= m_14_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1739 <= m_15_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1740 <= m_16_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1741 <= m_17_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1742 <= m_18_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1743 <= m_19_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1744 <= m_20_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1745 <= m_21_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1746 <= m_22_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1747 <= m_23_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1748 <= m_24_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1749 <= m_25_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1750 <= m_26_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1751 <= m_27_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1752 <= m_28_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1753 <= m_29_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1754 <= m_30_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1755 <= m_31_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1756 <= m_32_io_p[21]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1757 <= _T_796; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1758 <= m_11_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1759 <= m_12_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1760 <= m_13_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1761 <= m_14_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1762 <= m_15_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1763 <= m_16_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1764 <= m_17_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1765 <= m_18_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1766 <= m_19_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1767 <= m_20_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1768 <= m_21_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1769 <= m_22_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1770 <= m_23_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1771 <= m_24_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1772 <= m_25_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1773 <= m_26_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1774 <= m_27_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1775 <= m_28_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1776 <= m_29_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1777 <= m_30_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1778 <= m_31_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1779 <= m_32_io_p[22]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1781 <= m_11_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1782 <= m_12_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1783 <= m_13_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1784 <= m_14_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1785 <= m_15_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1786 <= m_16_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1787 <= m_17_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1788 <= m_18_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1789 <= m_19_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1790 <= m_20_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1791 <= m_21_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1792 <= m_22_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1793 <= m_23_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1794 <= m_24_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1795 <= m_25_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1796 <= m_26_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1797 <= m_27_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1798 <= m_28_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1799 <= m_29_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1800 <= m_30_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1801 <= m_31_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1802 <= m_32_io_p[23]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1803 <= _T_867; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1804 <= m_12_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1805 <= m_13_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1806 <= m_14_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1807 <= m_15_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1808 <= m_16_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1809 <= m_17_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1810 <= m_18_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1811 <= m_19_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1812 <= m_20_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1813 <= m_21_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1814 <= m_22_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1815 <= m_23_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1816 <= m_24_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1817 <= m_25_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1818 <= m_26_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1819 <= m_27_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1820 <= m_28_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1821 <= m_29_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1822 <= m_30_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1823 <= m_31_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1824 <= m_32_io_p[24]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1826 <= m_12_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1827 <= m_13_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1828 <= m_14_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1829 <= m_15_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1830 <= m_16_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1831 <= m_17_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1832 <= m_18_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1833 <= m_19_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1834 <= m_20_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1835 <= m_21_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1836 <= m_22_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1837 <= m_23_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1838 <= m_24_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1839 <= m_25_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1840 <= m_26_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1841 <= m_27_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1842 <= m_28_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1843 <= m_29_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1844 <= m_30_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1845 <= m_31_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1846 <= m_32_io_p[25]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1847 <= _T_938; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1848 <= m_13_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1849 <= m_14_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1850 <= m_15_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1851 <= m_16_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1852 <= m_17_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1853 <= m_18_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1854 <= m_19_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1855 <= m_20_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1856 <= m_21_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1857 <= m_22_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1858 <= m_23_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1859 <= m_24_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1860 <= m_25_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1861 <= m_26_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1862 <= m_27_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1863 <= m_28_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1864 <= m_29_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1865 <= m_30_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1866 <= m_31_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1867 <= m_32_io_p[26]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1869 <= m_13_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1870 <= m_14_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1871 <= m_15_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1872 <= m_16_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1873 <= m_17_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1874 <= m_18_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1875 <= m_19_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1876 <= m_20_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1877 <= m_21_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1878 <= m_22_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1879 <= m_23_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1880 <= m_24_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1881 <= m_25_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1882 <= m_26_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1883 <= m_27_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1884 <= m_28_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1885 <= m_29_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1886 <= m_30_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1887 <= m_31_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1888 <= m_32_io_p[27]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1889 <= _T_1009; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1890 <= m_14_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1891 <= m_15_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1892 <= m_16_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1893 <= m_17_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1894 <= m_18_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1895 <= m_19_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1896 <= m_20_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1897 <= m_21_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1898 <= m_22_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1899 <= m_23_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1900 <= m_24_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1901 <= m_25_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1902 <= m_26_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1903 <= m_27_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1904 <= m_28_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1905 <= m_29_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1906 <= m_30_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1907 <= m_31_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1908 <= m_32_io_p[28]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1910 <= m_14_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1911 <= m_15_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1912 <= m_16_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1913 <= m_17_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1914 <= m_18_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1915 <= m_19_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1916 <= m_20_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1917 <= m_21_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1918 <= m_22_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1919 <= m_23_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1920 <= m_24_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1921 <= m_25_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1922 <= m_26_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1923 <= m_27_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1924 <= m_28_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1925 <= m_29_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1926 <= m_30_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1927 <= m_31_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1928 <= m_32_io_p[29]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1929 <= _T_1080; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1930 <= m_15_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1931 <= m_16_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1932 <= m_17_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1933 <= m_18_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1934 <= m_19_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1935 <= m_20_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1936 <= m_21_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1937 <= m_22_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1938 <= m_23_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1939 <= m_24_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1940 <= m_25_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1941 <= m_26_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1942 <= m_27_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1943 <= m_28_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1944 <= m_29_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1945 <= m_30_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1946 <= m_31_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1947 <= m_32_io_p[30]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1949 <= m_15_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1950 <= m_16_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1951 <= m_17_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1952 <= m_18_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1953 <= m_19_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1954 <= m_20_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1955 <= m_21_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1956 <= m_22_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1957 <= m_23_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1958 <= m_24_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1959 <= m_25_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1960 <= m_26_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1961 <= m_27_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1962 <= m_28_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1963 <= m_29_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1964 <= m_30_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1965 <= m_31_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1966 <= m_32_io_p[31]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1967 <= _T_1151; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1968 <= m_16_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1969 <= m_17_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1970 <= m_18_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1971 <= m_19_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1972 <= m_20_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1973 <= m_21_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1974 <= m_22_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1975 <= m_23_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1976 <= m_24_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1977 <= m_25_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1978 <= m_26_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1979 <= m_27_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1980 <= m_28_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1981 <= m_29_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1982 <= m_30_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1983 <= m_31_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1984 <= m_32_io_p[32]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1986 <= m_16_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1987 <= m_17_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1988 <= m_18_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1989 <= m_19_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1990 <= m_20_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1991 <= m_21_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1992 <= m_22_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1993 <= m_23_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1994 <= m_24_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1995 <= m_25_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1996 <= m_26_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1997 <= m_27_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1998 <= m_28_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_1999 <= m_29_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2000 <= m_30_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2001 <= m_31_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2002 <= m_32_io_p[33]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2003 <= _T_1222; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2004 <= m_17_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2005 <= m_18_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2006 <= m_19_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2007 <= m_20_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2008 <= m_21_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2009 <= m_22_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2010 <= m_23_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2011 <= m_24_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2012 <= m_25_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2013 <= m_26_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2014 <= m_27_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2015 <= m_28_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2016 <= m_29_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2017 <= m_30_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2018 <= m_31_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2019 <= m_32_io_p[34]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2021 <= m_17_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2022 <= m_18_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2023 <= m_19_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2024 <= m_20_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2025 <= m_21_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2026 <= m_22_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2027 <= m_23_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2028 <= m_24_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2029 <= m_25_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2030 <= m_26_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2031 <= m_27_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2032 <= m_28_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2033 <= m_29_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2034 <= m_30_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2035 <= m_31_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2036 <= m_32_io_p[35]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2037 <= _T_1293; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2038 <= m_18_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2039 <= m_19_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2040 <= m_20_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2041 <= m_21_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2042 <= m_22_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2043 <= m_23_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2044 <= m_24_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2045 <= m_25_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2046 <= m_26_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2047 <= m_27_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2048 <= m_28_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2049 <= m_29_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2050 <= m_30_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2051 <= m_31_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2052 <= m_32_io_p[36]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2054 <= m_18_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2055 <= m_19_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2056 <= m_20_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2057 <= m_21_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2058 <= m_22_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2059 <= m_23_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2060 <= m_24_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2061 <= m_25_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2062 <= m_26_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2063 <= m_27_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2064 <= m_28_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2065 <= m_29_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2066 <= m_30_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2067 <= m_31_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2068 <= m_32_io_p[37]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2069 <= _T_1364; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2070 <= m_19_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2071 <= m_20_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2072 <= m_21_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2073 <= m_22_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2074 <= m_23_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2075 <= m_24_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2076 <= m_25_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2077 <= m_26_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2078 <= m_27_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2079 <= m_28_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2080 <= m_29_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2081 <= m_30_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2082 <= m_31_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2083 <= m_32_io_p[38]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2085 <= m_19_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2086 <= m_20_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2087 <= m_21_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2088 <= m_22_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2089 <= m_23_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2090 <= m_24_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2091 <= m_25_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2092 <= m_26_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2093 <= m_27_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2094 <= m_28_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2095 <= m_29_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2096 <= m_30_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2097 <= m_31_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2098 <= m_32_io_p[39]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2099 <= _T_1435; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2100 <= m_20_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2101 <= m_21_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2102 <= m_22_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2103 <= m_23_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2104 <= m_24_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2105 <= m_25_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2106 <= m_26_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2107 <= m_27_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2108 <= m_28_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2109 <= m_29_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2110 <= m_30_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2111 <= m_31_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2112 <= m_32_io_p[40]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2114 <= m_20_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2115 <= m_21_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2116 <= m_22_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2117 <= m_23_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2118 <= m_24_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2119 <= m_25_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2120 <= m_26_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2121 <= m_27_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2122 <= m_28_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2123 <= m_29_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2124 <= m_30_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2125 <= m_31_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2126 <= m_32_io_p[41]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2127 <= _T_1506; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2128 <= m_21_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2129 <= m_22_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2130 <= m_23_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2131 <= m_24_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2132 <= m_25_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2133 <= m_26_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2134 <= m_27_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2135 <= m_28_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2136 <= m_29_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2137 <= m_30_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2138 <= m_31_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2139 <= m_32_io_p[42]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2141 <= m_21_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2142 <= m_22_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2143 <= m_23_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2144 <= m_24_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2145 <= m_25_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2146 <= m_26_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2147 <= m_27_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2148 <= m_28_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2149 <= m_29_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2150 <= m_30_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2151 <= m_31_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2152 <= m_32_io_p[43]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2153 <= _T_1577; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2154 <= m_22_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2155 <= m_23_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2156 <= m_24_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2157 <= m_25_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2158 <= m_26_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2159 <= m_27_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2160 <= m_28_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2161 <= m_29_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2162 <= m_30_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2163 <= m_31_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2164 <= m_32_io_p[44]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2166 <= m_22_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2167 <= m_23_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2168 <= m_24_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2169 <= m_25_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2170 <= m_26_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2171 <= m_27_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2172 <= m_28_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2173 <= m_29_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2174 <= m_30_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2175 <= m_31_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2176 <= m_32_io_p[45]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2177 <= _T_1648; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2178 <= m_23_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2179 <= m_24_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2180 <= m_25_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2181 <= m_26_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2182 <= m_27_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2183 <= m_28_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2184 <= m_29_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2185 <= m_30_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2186 <= m_31_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2187 <= m_32_io_p[46]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2189 <= m_23_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2190 <= m_24_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2191 <= m_25_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2192 <= m_26_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2193 <= m_27_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2194 <= m_28_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2195 <= m_29_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2196 <= m_30_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2197 <= m_31_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2198 <= m_32_io_p[47]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2199 <= _T_1719; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2200 <= m_24_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2201 <= m_25_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2202 <= m_26_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2203 <= m_27_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2204 <= m_28_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2205 <= m_29_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2206 <= m_30_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2207 <= m_31_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2208 <= m_32_io_p[48]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2210 <= m_24_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2211 <= m_25_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2212 <= m_26_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2213 <= m_27_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2214 <= m_28_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2215 <= m_29_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2216 <= m_30_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2217 <= m_31_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2218 <= m_32_io_p[49]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2219 <= _T_1790; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2220 <= m_25_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2221 <= m_26_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2222 <= m_27_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2223 <= m_28_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2224 <= m_29_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2225 <= m_30_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2226 <= m_31_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2227 <= m_32_io_p[50]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2229 <= m_25_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2230 <= m_26_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2231 <= m_27_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2232 <= m_28_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2233 <= m_29_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2234 <= m_30_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2235 <= m_31_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2236 <= m_32_io_p[51]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2237 <= _T_1861; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2238 <= m_26_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2239 <= m_27_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2240 <= m_28_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2241 <= m_29_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2242 <= m_30_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2243 <= m_31_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2244 <= m_32_io_p[52]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2246 <= m_26_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2247 <= m_27_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2248 <= m_28_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2249 <= m_29_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2250 <= m_30_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2251 <= m_31_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2252 <= m_32_io_p[53]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2253 <= _T_1932; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2254 <= m_27_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2255 <= m_28_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2256 <= m_29_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2257 <= m_30_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2258 <= m_31_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2259 <= m_32_io_p[54]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2261 <= m_27_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2262 <= m_28_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2263 <= m_29_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2264 <= m_30_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2265 <= m_31_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2266 <= m_32_io_p[55]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2267 <= _T_2003; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2268 <= m_28_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2269 <= m_29_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2270 <= m_30_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2271 <= m_31_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2272 <= m_32_io_p[56]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2274 <= m_28_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2275 <= m_29_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2276 <= m_30_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2277 <= m_31_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2278 <= m_32_io_p[57]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2279 <= _T_2074; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2280 <= m_29_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2281 <= m_30_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2282 <= m_31_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2283 <= m_32_io_p[58]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2285 <= m_29_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2286 <= m_30_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2287 <= m_31_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2288 <= m_32_io_p[59]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2289 <= _T_2145; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2290 <= m_30_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2291 <= m_31_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2292 <= m_32_io_p[60]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2294 <= m_30_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2295 <= m_31_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2296 <= m_32_io_p[61]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2297 <= _T_2216; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2298 <= m_31_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2299 <= m_32_io_p[62]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2301 <= m_31_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2302 <= m_32_io_p[63]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2303 <= _T_2287; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2304 <= m_32_io_p[64]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2306 <= m_32_io_p[65]; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2307 <= _T_2358; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2308 <= m_33_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2309 <= m_803_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2310 <= m_1329_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2311 <= m_1698_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2312 <= m_1699_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2313 <= m_1698_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2314 <= m_1700_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2315 <= m_1699_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2316 <= m_1701_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2317 <= m_1700_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2318 <= m_1702_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2319 <= m_1701_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2320 <= m_1703_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2321 <= m_1702_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2322 <= m_1704_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2323 <= m_1703_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2324 <= m_1705_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2325 <= m_1704_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2326 <= s_0_366; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2327 <= m_1705_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2328 <= s_0_367; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2329 <= c_0_366; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2330 <= s_0_368; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2331 <= c_0_367; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2332 <= s_0_369; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2333 <= c_0_368; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2334 <= s_0_370; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2335 <= c_0_369; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2336 <= s_0_371; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2337 <= c_0_370; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2338 <= s_0_372; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2339 <= c_0_371; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2340 <= m_1344_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2341 <= s_0_373; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2342 <= c_0_372; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2343 <= m_1346_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2344 <= s_0_374; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2345 <= c_0_373; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2346 <= m_1348_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2347 <= s_0_375; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2348 <= c_0_374; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2349 <= m_1350_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2350 <= s_0_376; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2351 <= c_0_375; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2352 <= c_1_220; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2353 <= s_0_377; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2354 <= c_0_376; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2355 <= c_1_221; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2356 <= s_0_378; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2357 <= c_0_377; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2358 <= c_1_222; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2359 <= s_0_379; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2360 <= c_0_378; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2361 <= c_1_223; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2362 <= s_0_380; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2363 <= c_0_379; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2364 <= m_1721_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2365 <= s_0_381; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2366 <= c_0_380; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2367 <= m_1723_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2368 <= m_1721_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2369 <= s_0_382; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2370 <= c_0_381; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2371 <= m_1725_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2372 <= m_1723_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2373 <= s_0_383; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2374 <= c_0_382; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2375 <= m_1727_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2376 <= m_1725_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2377 <= s_0_384; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2378 <= c_0_383; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2379 <= m_1729_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2380 <= m_1727_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2381 <= s_0_385; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2382 <= c_0_384; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2383 <= s_2_314; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2384 <= m_1729_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2385 <= s_0_386; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2386 <= c_0_385; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2387 <= s_2_315; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2388 <= c_1_314; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2389 <= s_0_387; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2390 <= c_0_386; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2391 <= s_2_316; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2392 <= c_1_315; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2393 <= s_0_388; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2394 <= c_0_387; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2395 <= s_2_317; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2396 <= c_1_316; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2397 <= s_0_389; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2398 <= c_0_388; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2399 <= s_2_318; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2400 <= c_1_317; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2401 <= s_0_390; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2402 <= c_0_389; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2403 <= s_2_319; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2404 <= c_1_318; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2405 <= s_0_391; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2406 <= c_0_390; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2407 <= s_2_320; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2408 <= c_1_319; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2409 <= s_0_392; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2410 <= c_0_391; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2411 <= s_2_321; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2412 <= c_1_320; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2413 <= s_0_393; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2414 <= c_0_392; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2415 <= s_2_322; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2416 <= c_1_321; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2417 <= m_897_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2418 <= s_0_394; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2419 <= c_0_393; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2420 <= s_2_323; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2421 <= c_1_322; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2422 <= m_902_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2423 <= s_0_395; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2424 <= c_0_394; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2425 <= s_2_324; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2426 <= c_1_323; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2427 <= m_907_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2428 <= s_0_396; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2429 <= c_0_395; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2430 <= s_2_325; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2431 <= c_1_324; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2432 <= c_4_78; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2433 <= s_0_397; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2434 <= c_0_396; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2435 <= s_2_326; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2436 <= c_1_325; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2437 <= c_4_79; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2438 <= s_0_398; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2439 <= c_0_397; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2440 <= s_2_327; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2441 <= c_1_326; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2442 <= m_1414_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2443 <= s_0_399; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2444 <= c_0_398; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2445 <= s_2_328; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2446 <= c_1_327; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2447 <= m_1760_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2448 <= s_0_400; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2449 <= c_0_399; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2450 <= s_2_329; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2451 <= c_1_328; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2452 <= m_1763_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2453 <= m_1760_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2454 <= s_0_401; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2455 <= c_0_400; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2456 <= s_2_330; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2457 <= c_1_329; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2458 <= m_1766_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2459 <= m_1763_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2460 <= s_0_402; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2461 <= c_0_401; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2462 <= s_2_331; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2463 <= c_1_330; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2464 <= m_1769_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2465 <= m_1766_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2466 <= s_0_403; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2467 <= c_0_402; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2468 <= s_2_332; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2469 <= c_1_331; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2470 <= m_1772_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2471 <= m_1769_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2472 <= s_0_404; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2473 <= c_0_403; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2474 <= s_2_333; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2475 <= c_1_332; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2476 <= m_1775_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2477 <= m_1772_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2478 <= s_0_405; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2479 <= c_0_404; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2480 <= s_2_334; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2481 <= c_1_333; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2482 <= m_1778_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2483 <= m_1775_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2484 <= s_0_406; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2485 <= c_0_405; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2486 <= s_2_335; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2487 <= c_1_334; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2488 <= m_1781_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2489 <= m_1778_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2490 <= s_0_407; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2491 <= c_0_406; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2492 <= s_2_336; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2493 <= c_1_335; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2494 <= s_4_250; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2495 <= m_1781_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2496 <= s_0_408; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2497 <= c_0_407; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2498 <= s_2_337; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2499 <= c_1_336; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2500 <= s_4_251; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2501 <= c_2_250; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2502 <= s_0_409; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2503 <= c_0_408; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2504 <= s_2_338; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2505 <= c_1_337; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2506 <= s_4_252; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2507 <= c_2_251; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2508 <= s_0_410; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2509 <= c_0_409; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2510 <= s_2_339; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2511 <= c_1_338; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2512 <= s_4_253; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2513 <= c_2_252; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2514 <= s_0_411; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2515 <= c_0_410; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2516 <= s_2_340; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2517 <= c_1_339; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2518 <= s_4_254; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2519 <= c_2_253; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2520 <= s_0_412; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2521 <= c_0_411; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2522 <= s_2_341; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2523 <= c_1_340; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2524 <= s_4_255; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2525 <= c_2_254; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2526 <= m_1467_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2527 <= s_0_413; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2528 <= c_0_412; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2529 <= s_2_342; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2530 <= c_1_341; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2531 <= s_4_256; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2532 <= c_2_255; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2533 <= m_1472_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2534 <= s_0_414; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2535 <= c_0_413; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2536 <= s_2_343; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2537 <= c_1_342; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2538 <= s_4_257; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2539 <= c_2_256; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2540 <= m_1477_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2541 <= s_0_415; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2542 <= c_0_414; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2543 <= s_2_344; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2544 <= c_1_343; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2545 <= s_4_258; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2546 <= c_2_257; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2547 <= m_1482_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2548 <= s_0_416; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2549 <= c_0_415; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2550 <= s_2_345; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2551 <= c_1_344; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2552 <= s_4_259; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2553 <= c_2_258; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2554 <= m_1487_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2555 <= s_0_417; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2556 <= c_0_416; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2557 <= s_2_346; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2558 <= c_1_345; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2559 <= s_4_260; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2560 <= c_2_259; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2561 <= c_4_128; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2562 <= s_0_418; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2563 <= c_0_417; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2564 <= s_2_347; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2565 <= c_1_346; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2566 <= s_4_261; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2567 <= c_2_260; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2568 <= c_4_129; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2569 <= s_0_419; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2570 <= c_0_418; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2571 <= s_2_348; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2572 <= c_1_347; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2573 <= s_4_262; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2574 <= c_2_261; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2575 <= c_4_130; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2576 <= s_0_420; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2577 <= c_0_419; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2578 <= s_2_349; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2579 <= c_1_348; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2580 <= s_4_263; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2581 <= c_2_262; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2582 <= c_4_131; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2583 <= s_0_421; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2584 <= c_0_420; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2585 <= s_2_350; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2586 <= c_1_349; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2587 <= s_4_264; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2588 <= c_2_263; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2589 <= c_4_132; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2590 <= s_0_422; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2591 <= c_0_421; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2592 <= s_2_351; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2593 <= c_1_350; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2594 <= s_4_265; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2595 <= c_2_264; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2596 <= c_4_133; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2597 <= s_0_423; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2598 <= c_0_422; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2599 <= s_2_352; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2600 <= c_1_351; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2601 <= s_4_266; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2602 <= c_2_265; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2603 <= c_4_134; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2604 <= s_0_424; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2605 <= c_0_423; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2606 <= s_2_353; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2607 <= c_1_352; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2608 <= s_4_267; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2609 <= c_2_266; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2610 <= c_4_135; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2611 <= s_0_425; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2612 <= c_0_424; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2613 <= s_2_354; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2614 <= c_1_353; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2615 <= s_4_268; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2616 <= c_2_267; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2617 <= c_4_136; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2618 <= s_0_426; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2619 <= c_0_425; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2620 <= s_2_355; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2621 <= c_1_354; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2622 <= s_4_269; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2623 <= c_2_268; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2624 <= c_4_137; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2625 <= s_0_427; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2626 <= c_0_426; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2627 <= s_2_356; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2628 <= c_1_355; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2629 <= s_4_270; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2630 <= c_2_269; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2631 <= m_1542_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2632 <= s_0_428; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2633 <= c_0_427; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2634 <= s_2_357; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2635 <= c_1_356; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2636 <= s_4_271; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2637 <= c_2_270; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2638 <= m_1547_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2639 <= s_0_429; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2640 <= c_0_428; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2641 <= s_2_358; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2642 <= c_1_357; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2643 <= s_4_272; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2644 <= c_2_271; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2645 <= m_1552_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2646 <= s_0_430; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2647 <= c_0_429; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2648 <= s_2_359; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2649 <= c_1_358; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2650 <= s_4_273; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2651 <= c_2_272; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2652 <= m_1557_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2653 <= s_0_431; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2654 <= c_0_430; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2655 <= s_2_360; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2656 <= c_1_359; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2657 <= s_4_274; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2658 <= c_2_273; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2659 <= m_1562_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2660 <= s_0_432; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2661 <= c_0_431; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2662 <= s_2_361; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2663 <= c_1_360; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2664 <= s_4_275; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2665 <= c_2_274; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2666 <= m_1567_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2667 <= s_0_433; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2668 <= c_0_432; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2669 <= s_2_362; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2670 <= c_1_361; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2671 <= s_4_276; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2672 <= c_2_275; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2673 <= s_0_434; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2674 <= c_0_433; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2675 <= s_2_363; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2676 <= c_1_362; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2677 <= m_1865_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2678 <= c_2_276; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2679 <= s_0_435; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2680 <= c_0_434; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2681 <= s_2_364; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2682 <= c_1_363; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2683 <= m_1868_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2684 <= m_1865_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2685 <= s_0_436; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2686 <= c_0_435; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2687 <= s_2_365; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2688 <= c_1_364; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2689 <= m_1871_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2690 <= m_1868_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2691 <= s_0_437; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2692 <= c_0_436; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2693 <= s_2_366; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2694 <= c_1_365; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2695 <= m_1874_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2696 <= m_1871_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2697 <= s_0_438; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2698 <= c_0_437; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2699 <= s_2_367; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2700 <= c_1_366; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2701 <= m_1877_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2702 <= m_1874_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2703 <= s_0_439; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2704 <= c_0_438; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2705 <= s_2_368; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2706 <= c_1_367; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2707 <= m_1880_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2708 <= m_1877_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2709 <= s_0_440; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2710 <= c_0_439; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2711 <= s_2_369; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2712 <= c_1_368; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2713 <= m_1883_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2714 <= m_1880_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2715 <= s_0_441; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2716 <= c_0_440; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2717 <= s_2_370; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2718 <= c_1_369; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2719 <= m_1886_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2720 <= m_1883_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2721 <= s_0_442; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2722 <= c_0_441; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2723 <= s_2_371; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2724 <= c_1_370; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2725 <= m_1889_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2726 <= m_1886_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2727 <= s_0_443; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2728 <= c_0_442; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2729 <= s_2_372; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2730 <= c_1_371; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2731 <= m_1892_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2732 <= m_1889_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2733 <= s_0_444; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2734 <= c_0_443; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2735 <= s_2_373; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2736 <= c_1_372; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2737 <= m_1895_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2738 <= m_1892_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2739 <= s_0_445; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2740 <= c_0_444; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2741 <= s_2_374; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2742 <= c_1_373; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2743 <= c_4_127; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2744 <= m_1895_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2745 <= s_0_446; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2746 <= c_0_445; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2747 <= s_2_375; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2748 <= c_1_374; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2749 <= m_1222_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2750 <= s_0_447; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2751 <= c_0_446; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2752 <= s_2_376; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2753 <= c_1_375; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2754 <= m_1227_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2755 <= s_0_448; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2756 <= c_0_447; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2757 <= s_2_377; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2758 <= c_1_376; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2759 <= m_1232_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2760 <= s_0_449; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2761 <= c_0_448; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2762 <= s_2_378; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2763 <= c_1_377; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2764 <= m_1237_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2765 <= s_0_450; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2766 <= c_0_449; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2767 <= s_2_379; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2768 <= c_1_378; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2769 <= m_1242_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2770 <= s_0_451; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2771 <= c_0_450; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2772 <= s_2_380; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2773 <= c_1_379; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2774 <= s_0_452; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2775 <= c_0_451; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2776 <= s_2_381; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2777 <= c_1_380; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2778 <= s_0_453; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2779 <= c_0_452; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2780 <= s_2_382; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2781 <= c_1_381; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2782 <= s_0_454; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2783 <= c_0_453; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2784 <= s_2_383; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2785 <= c_1_382; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2786 <= s_0_455; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2787 <= c_0_454; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2788 <= s_2_384; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2789 <= c_1_383; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2790 <= s_0_456; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2791 <= c_0_455; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2792 <= s_2_385; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2793 <= c_1_384; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2794 <= s_0_457; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2795 <= c_0_456; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2796 <= s_2_386; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2797 <= c_1_385; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2798 <= s_0_458; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2799 <= c_0_457; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2800 <= s_2_387; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2801 <= c_1_386; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2802 <= s_0_459; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2803 <= c_0_458; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2804 <= m_1925_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2805 <= c_1_387; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2806 <= s_0_460; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2807 <= c_0_459; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2808 <= m_1927_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2809 <= m_1925_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2810 <= s_0_461; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2811 <= c_0_460; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2812 <= m_1929_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2813 <= m_1927_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2814 <= s_0_462; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2815 <= c_0_461; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2816 <= c_1_306; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2817 <= m_1929_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2818 <= s_0_463; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2819 <= c_0_462; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2820 <= c_1_307; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2821 <= s_0_464; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2822 <= c_0_463; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2823 <= c_1_308; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2824 <= s_0_465; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2825 <= c_0_464; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2826 <= c_1_309; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2827 <= s_0_466; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2828 <= c_0_465; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2829 <= c_1_310; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2830 <= s_0_467; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2831 <= c_0_466; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2832 <= c_1_311; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2833 <= s_0_468; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2834 <= c_0_467; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2835 <= c_1_312; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2836 <= s_0_469; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2837 <= c_0_468; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2838 <= c_1_313; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2839 <= s_0_470; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2840 <= c_0_469; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2841 <= s_0_471; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2842 <= c_0_470; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2843 <= s_0_472; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2844 <= c_0_471; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2845 <= s_0_473; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2846 <= c_0_472; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2847 <= s_0_474; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2848 <= c_0_473; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2849 <= s_0_475; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2850 <= c_0_474; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2851 <= m_1944_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2852 <= c_0_475; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2853 <= m_1945_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2854 <= m_1944_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2855 <= m_1946_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2856 <= m_1945_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2857 <= m_1947_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2858 <= m_1946_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2859 <= m_1948_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2860 <= m_1947_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2861 <= m_1949_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2862 <= m_1948_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2863 <= m_1950_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2864 <= m_1949_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2865 <= m_1951_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2866 <= m_1950_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2867 <= m_1952_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2868 <= m_1951_io_out_1; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2869 <= m_1953_io_out_0; // @[Reg.scala 17:22]
    end
    if (io_in_valid) begin // @[Reg.scala 17:18]
      r_2870 <= m_1952_io_out_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[MUL.scala 334:22]
      count <= 8'h0; // @[MUL.scala 334:22]
    end else if (io_in_valid & ~io_out_valid) begin // @[MUL.scala 336:15]
      count <= _count_T_5;
    end else begin
      count <= 8'h0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  r_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  r_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  r_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  r_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  r_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  r_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  r_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  r_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  r_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  r_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  r_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  r_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  r_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  r_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  r_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  r_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  r_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  r_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  r_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  r_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  r_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  r_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  r_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  r_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  r_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  r_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  r_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  r_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  r_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  r_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  r_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  r_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  r_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  r_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  r_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  r_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  r_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  r_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  r_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  r_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  r_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  r_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  r_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  r_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  r_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  r_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  r_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  r_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  r_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  r_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  r_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  r_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  r_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  r_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  r_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  r_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  r_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  r_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  r_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  r_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  r_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  r_63 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  r_64 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  r_65 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  r_66 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  r_67 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  r_68 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  r_69 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  r_70 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  r_71 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  r_72 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  r_73 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  r_74 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  r_75 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  r_76 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  r_77 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  r_78 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  r_79 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  r_80 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  r_81 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  r_82 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  r_83 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  r_84 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  r_85 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  r_86 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  r_87 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  r_88 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  r_89 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  r_90 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  r_91 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  r_92 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  r_93 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  r_94 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  r_95 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  r_96 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  r_97 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  r_98 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  r_99 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  r_100 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  r_101 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  r_102 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  r_103 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  r_104 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  r_105 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  r_106 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  r_107 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  r_108 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  r_109 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  r_110 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  r_111 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  r_112 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  r_113 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  r_114 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  r_115 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  r_116 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  r_117 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  r_118 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  r_119 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  r_120 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  r_121 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  r_122 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  r_123 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  r_124 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  r_125 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  r_126 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  r_127 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  r_128 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  r_129 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  r_130 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  r_131 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  r_132 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  r_133 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  r_134 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  r_135 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  r_136 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  r_137 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  r_138 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  r_139 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  r_140 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  r_141 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  r_142 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  r_143 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  r_144 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  r_145 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  r_146 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  r_147 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  r_148 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  r_149 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  r_150 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  r_151 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  r_152 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  r_153 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  r_154 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  r_155 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  r_156 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  r_157 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  r_158 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  r_159 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  r_160 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  r_161 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  r_162 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  r_163 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  r_164 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  r_165 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  r_166 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  r_167 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  r_168 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  r_169 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  r_170 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  r_171 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  r_172 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  r_173 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  r_174 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  r_175 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  r_176 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  r_177 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  r_178 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  r_179 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  r_180 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  r_181 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  r_182 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  r_183 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  r_184 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  r_185 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  r_186 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  r_187 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  r_188 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  r_189 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  r_190 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  r_191 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  r_192 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  r_193 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  r_194 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  r_195 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  r_196 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  r_197 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  r_198 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  r_199 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  r_200 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  r_201 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  r_202 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  r_203 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  r_204 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  r_205 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  r_206 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  r_207 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  r_208 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  r_209 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  r_210 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  r_211 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  r_212 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  r_213 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  r_214 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  r_215 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  r_216 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  r_217 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  r_218 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  r_219 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  r_220 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  r_221 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  r_222 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  r_223 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  r_224 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  r_225 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  r_226 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  r_227 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  r_228 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  r_229 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  r_230 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  r_231 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  r_232 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  r_233 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  r_234 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  r_235 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  r_236 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  r_237 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  r_238 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  r_239 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  r_240 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  r_241 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  r_242 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  r_243 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  r_244 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  r_245 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  r_246 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  r_247 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  r_248 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  r_249 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  r_250 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  r_251 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  r_252 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  r_253 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  r_254 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  r_255 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  r_256 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  r_257 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  r_258 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  r_259 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  r_260 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  r_261 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  r_262 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  r_263 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  r_264 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  r_265 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  r_266 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  r_267 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  r_268 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  r_269 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  r_270 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  r_271 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  r_272 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  r_273 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  r_274 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  r_275 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  r_276 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  r_277 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  r_278 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  r_279 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  r_280 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  r_281 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  r_282 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  r_283 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  r_284 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  r_285 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  r_286 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  r_287 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  r_288 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  r_289 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  r_290 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  r_291 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  r_292 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  r_293 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  r_294 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  r_295 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  r_296 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  r_297 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  r_298 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  r_299 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  r_300 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  r_301 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  r_302 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  r_303 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  r_304 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  r_305 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  r_306 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  r_307 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  r_308 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  r_309 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  r_310 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  r_311 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  r_312 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  r_313 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  r_314 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  r_315 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  r_316 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  r_317 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  r_318 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  r_319 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  r_320 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  r_321 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  r_322 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  r_323 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  r_324 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  r_325 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  r_326 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  r_327 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  r_328 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  r_329 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  r_330 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  r_331 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  r_332 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  r_333 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  r_334 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  r_335 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  r_336 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  r_337 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  r_338 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  r_339 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  r_340 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  r_341 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  r_342 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  r_343 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  r_344 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  r_345 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  r_346 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  r_347 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  r_348 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  r_349 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  r_350 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  r_351 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  r_352 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  r_353 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  r_354 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  r_355 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  r_356 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  r_357 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  r_358 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  r_359 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  r_360 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  r_361 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  r_362 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  r_363 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  r_364 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  r_365 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  r_366 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  r_367 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  r_368 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  r_369 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  r_370 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  r_371 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  r_372 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  r_373 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  r_374 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  r_375 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  r_376 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  r_377 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  r_378 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  r_379 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  r_380 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  r_381 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  r_382 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  r_383 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  r_384 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  r_385 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  r_386 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  r_387 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  r_388 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  r_389 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  r_390 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  r_391 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  r_392 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  r_393 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  r_394 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  r_395 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  r_396 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  r_397 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  r_398 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  r_399 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  r_400 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  r_401 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  r_402 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  r_403 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  r_404 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  r_405 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  r_406 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  r_407 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  r_408 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  r_409 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  r_410 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  r_411 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  r_412 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  r_413 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  r_414 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  r_415 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  r_416 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  r_417 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  r_418 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  r_419 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  r_420 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  r_421 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  r_422 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  r_423 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  r_424 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  r_425 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  r_426 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  r_427 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  r_428 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  r_429 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  r_430 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  r_431 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  r_432 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  r_433 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  r_434 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  r_435 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  r_436 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  r_437 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  r_438 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  r_439 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  r_440 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  r_441 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  r_442 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  r_443 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  r_444 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  r_445 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  r_446 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  r_447 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  r_448 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  r_449 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  r_450 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  r_451 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  r_452 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  r_453 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  r_454 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  r_455 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  r_456 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  r_457 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  r_458 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  r_459 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  r_460 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  r_461 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  r_462 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  r_463 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  r_464 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  r_465 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  r_466 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  r_467 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  r_468 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  r_469 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  r_470 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  r_471 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  r_472 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  r_473 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  r_474 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  r_475 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  r_476 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  r_477 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  r_478 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  r_479 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  r_480 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  r_481 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  r_482 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  r_483 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  r_484 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  r_485 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  r_486 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  r_487 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  r_488 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  r_489 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  r_490 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  r_491 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  r_492 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  r_493 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  r_494 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  r_495 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  r_496 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  r_497 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  r_498 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  r_499 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  r_500 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  r_501 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  r_502 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  r_503 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  r_504 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  r_505 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  r_506 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  r_507 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  r_508 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  r_509 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  r_510 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  r_511 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  r_512 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  r_513 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  r_514 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  r_515 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  r_516 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  r_517 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  r_518 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  r_519 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  r_520 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  r_521 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  r_522 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  r_523 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  r_524 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  r_525 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  r_526 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  r_527 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  r_528 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  r_529 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  r_530 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  r_531 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  r_532 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  r_533 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  r_534 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  r_535 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  r_536 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  r_537 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  r_538 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  r_539 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  r_540 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  r_541 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  r_542 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  r_543 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  r_544 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  r_545 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  r_546 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  r_547 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  r_548 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  r_549 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  r_550 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  r_551 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  r_552 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  r_553 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  r_554 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  r_555 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  r_556 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  r_557 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  r_558 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  r_559 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  r_560 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  r_561 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  r_562 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  r_563 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  r_564 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  r_565 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  r_566 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  r_567 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  r_568 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  r_569 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  r_570 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  r_571 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  r_572 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  r_573 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  r_574 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  r_575 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  r_576 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  r_577 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  r_578 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  r_579 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  r_580 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  r_581 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  r_582 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  r_583 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  r_584 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  r_585 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  r_586 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  r_587 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  r_588 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  r_589 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  r_590 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  r_591 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  r_592 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  r_593 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  r_594 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  r_595 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  r_596 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  r_597 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  r_598 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  r_599 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  r_600 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  r_601 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  r_602 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  r_603 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  r_604 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  r_605 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  r_606 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  r_607 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  r_608 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  r_609 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  r_610 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  r_611 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  r_612 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  r_613 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  r_614 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  r_615 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  r_616 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  r_617 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  r_618 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  r_619 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  r_620 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  r_621 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  r_622 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  r_623 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  r_624 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  r_625 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  r_626 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  r_627 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  r_628 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  r_629 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  r_630 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  r_631 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  r_632 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  r_633 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  r_634 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  r_635 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  r_636 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  r_637 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  r_638 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  r_639 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  r_640 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  r_641 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  r_642 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  r_643 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  r_644 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  r_645 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  r_646 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  r_647 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  r_648 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  r_649 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  r_650 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  r_651 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  r_652 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  r_653 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  r_654 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  r_655 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  r_656 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  r_657 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  r_658 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  r_659 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  r_660 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  r_661 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  r_662 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  r_663 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  r_664 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  r_665 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  r_666 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  r_667 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  r_668 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  r_669 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  r_670 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  r_671 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  r_672 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  r_673 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  r_674 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  r_675 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  r_676 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  r_677 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  r_678 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  r_679 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  r_680 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  r_681 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  r_682 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  r_683 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  r_684 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  r_685 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  r_686 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  r_687 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  r_688 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  r_689 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  r_690 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  r_691 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  r_692 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  r_693 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  r_694 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  r_695 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  r_696 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  r_697 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  r_698 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  r_699 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  r_700 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  r_701 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  r_702 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  r_703 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  r_704 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  r_705 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  r_706 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  r_707 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  r_708 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  r_709 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  r_710 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  r_711 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  r_712 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  r_713 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  r_714 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  r_715 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  r_716 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  r_717 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  r_718 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  r_719 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  r_720 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  r_721 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  r_722 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  r_723 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  r_724 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  r_725 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  r_726 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  r_727 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  r_728 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  r_729 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  r_730 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  r_731 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  r_732 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  r_733 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  r_734 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  r_735 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  r_736 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  r_737 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  r_738 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  r_739 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  r_740 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  r_741 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  r_742 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  r_743 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  r_744 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  r_745 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  r_746 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  r_747 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  r_748 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  r_749 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  r_750 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  r_751 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  r_752 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  r_753 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  r_754 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  r_755 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  r_756 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  r_757 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  r_758 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  r_759 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  r_760 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  r_761 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  r_762 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  r_763 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  r_764 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  r_765 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  r_766 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  r_767 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  r_768 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  r_769 = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  r_770 = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  r_771 = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  r_772 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  r_773 = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  r_774 = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  r_775 = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  r_776 = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  r_777 = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  r_778 = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  r_779 = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  r_780 = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  r_781 = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  r_782 = _RAND_782[0:0];
  _RAND_783 = {1{`RANDOM}};
  r_783 = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  r_784 = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  r_785 = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  r_786 = _RAND_786[0:0];
  _RAND_787 = {1{`RANDOM}};
  r_787 = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  r_788 = _RAND_788[0:0];
  _RAND_789 = {1{`RANDOM}};
  r_789 = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  r_790 = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  r_791 = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  r_792 = _RAND_792[0:0];
  _RAND_793 = {1{`RANDOM}};
  r_793 = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  r_794 = _RAND_794[0:0];
  _RAND_795 = {1{`RANDOM}};
  r_795 = _RAND_795[0:0];
  _RAND_796 = {1{`RANDOM}};
  r_796 = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  r_797 = _RAND_797[0:0];
  _RAND_798 = {1{`RANDOM}};
  r_798 = _RAND_798[0:0];
  _RAND_799 = {1{`RANDOM}};
  r_799 = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  r_800 = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  r_801 = _RAND_801[0:0];
  _RAND_802 = {1{`RANDOM}};
  r_802 = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  r_803 = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  r_804 = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  r_805 = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  r_806 = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  r_807 = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  r_808 = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  r_809 = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  r_810 = _RAND_810[0:0];
  _RAND_811 = {1{`RANDOM}};
  r_811 = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  r_812 = _RAND_812[0:0];
  _RAND_813 = {1{`RANDOM}};
  r_813 = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  r_814 = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  r_815 = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  r_816 = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  r_817 = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  r_818 = _RAND_818[0:0];
  _RAND_819 = {1{`RANDOM}};
  r_819 = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  r_820 = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  r_821 = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  r_822 = _RAND_822[0:0];
  _RAND_823 = {1{`RANDOM}};
  r_823 = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  r_824 = _RAND_824[0:0];
  _RAND_825 = {1{`RANDOM}};
  r_825 = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  r_826 = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  r_827 = _RAND_827[0:0];
  _RAND_828 = {1{`RANDOM}};
  r_828 = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  r_829 = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  r_830 = _RAND_830[0:0];
  _RAND_831 = {1{`RANDOM}};
  r_831 = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  r_832 = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  r_833 = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  r_834 = _RAND_834[0:0];
  _RAND_835 = {1{`RANDOM}};
  r_835 = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  r_836 = _RAND_836[0:0];
  _RAND_837 = {1{`RANDOM}};
  r_837 = _RAND_837[0:0];
  _RAND_838 = {1{`RANDOM}};
  r_838 = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  r_839 = _RAND_839[0:0];
  _RAND_840 = {1{`RANDOM}};
  r_840 = _RAND_840[0:0];
  _RAND_841 = {1{`RANDOM}};
  r_841 = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  r_842 = _RAND_842[0:0];
  _RAND_843 = {1{`RANDOM}};
  r_843 = _RAND_843[0:0];
  _RAND_844 = {1{`RANDOM}};
  r_844 = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  r_845 = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  r_846 = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  r_847 = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  r_848 = _RAND_848[0:0];
  _RAND_849 = {1{`RANDOM}};
  r_849 = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  r_850 = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  r_851 = _RAND_851[0:0];
  _RAND_852 = {1{`RANDOM}};
  r_852 = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  r_853 = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  r_854 = _RAND_854[0:0];
  _RAND_855 = {1{`RANDOM}};
  r_855 = _RAND_855[0:0];
  _RAND_856 = {1{`RANDOM}};
  r_856 = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  r_857 = _RAND_857[0:0];
  _RAND_858 = {1{`RANDOM}};
  r_858 = _RAND_858[0:0];
  _RAND_859 = {1{`RANDOM}};
  r_859 = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  r_860 = _RAND_860[0:0];
  _RAND_861 = {1{`RANDOM}};
  r_861 = _RAND_861[0:0];
  _RAND_862 = {1{`RANDOM}};
  r_862 = _RAND_862[0:0];
  _RAND_863 = {1{`RANDOM}};
  r_863 = _RAND_863[0:0];
  _RAND_864 = {1{`RANDOM}};
  r_864 = _RAND_864[0:0];
  _RAND_865 = {1{`RANDOM}};
  r_865 = _RAND_865[0:0];
  _RAND_866 = {1{`RANDOM}};
  r_866 = _RAND_866[0:0];
  _RAND_867 = {1{`RANDOM}};
  r_867 = _RAND_867[0:0];
  _RAND_868 = {1{`RANDOM}};
  r_868 = _RAND_868[0:0];
  _RAND_869 = {1{`RANDOM}};
  r_869 = _RAND_869[0:0];
  _RAND_870 = {1{`RANDOM}};
  r_870 = _RAND_870[0:0];
  _RAND_871 = {1{`RANDOM}};
  r_871 = _RAND_871[0:0];
  _RAND_872 = {1{`RANDOM}};
  r_872 = _RAND_872[0:0];
  _RAND_873 = {1{`RANDOM}};
  r_873 = _RAND_873[0:0];
  _RAND_874 = {1{`RANDOM}};
  r_874 = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  r_875 = _RAND_875[0:0];
  _RAND_876 = {1{`RANDOM}};
  r_876 = _RAND_876[0:0];
  _RAND_877 = {1{`RANDOM}};
  r_877 = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  r_878 = _RAND_878[0:0];
  _RAND_879 = {1{`RANDOM}};
  r_879 = _RAND_879[0:0];
  _RAND_880 = {1{`RANDOM}};
  r_880 = _RAND_880[0:0];
  _RAND_881 = {1{`RANDOM}};
  r_881 = _RAND_881[0:0];
  _RAND_882 = {1{`RANDOM}};
  r_882 = _RAND_882[0:0];
  _RAND_883 = {1{`RANDOM}};
  r_883 = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  r_884 = _RAND_884[0:0];
  _RAND_885 = {1{`RANDOM}};
  r_885 = _RAND_885[0:0];
  _RAND_886 = {1{`RANDOM}};
  r_886 = _RAND_886[0:0];
  _RAND_887 = {1{`RANDOM}};
  r_887 = _RAND_887[0:0];
  _RAND_888 = {1{`RANDOM}};
  r_888 = _RAND_888[0:0];
  _RAND_889 = {1{`RANDOM}};
  r_889 = _RAND_889[0:0];
  _RAND_890 = {1{`RANDOM}};
  r_890 = _RAND_890[0:0];
  _RAND_891 = {1{`RANDOM}};
  r_891 = _RAND_891[0:0];
  _RAND_892 = {1{`RANDOM}};
  r_892 = _RAND_892[0:0];
  _RAND_893 = {1{`RANDOM}};
  r_893 = _RAND_893[0:0];
  _RAND_894 = {1{`RANDOM}};
  r_894 = _RAND_894[0:0];
  _RAND_895 = {1{`RANDOM}};
  r_895 = _RAND_895[0:0];
  _RAND_896 = {1{`RANDOM}};
  r_896 = _RAND_896[0:0];
  _RAND_897 = {1{`RANDOM}};
  r_897 = _RAND_897[0:0];
  _RAND_898 = {1{`RANDOM}};
  r_898 = _RAND_898[0:0];
  _RAND_899 = {1{`RANDOM}};
  r_899 = _RAND_899[0:0];
  _RAND_900 = {1{`RANDOM}};
  r_900 = _RAND_900[0:0];
  _RAND_901 = {1{`RANDOM}};
  r_901 = _RAND_901[0:0];
  _RAND_902 = {1{`RANDOM}};
  r_902 = _RAND_902[0:0];
  _RAND_903 = {1{`RANDOM}};
  r_903 = _RAND_903[0:0];
  _RAND_904 = {1{`RANDOM}};
  r_904 = _RAND_904[0:0];
  _RAND_905 = {1{`RANDOM}};
  r_905 = _RAND_905[0:0];
  _RAND_906 = {1{`RANDOM}};
  r_906 = _RAND_906[0:0];
  _RAND_907 = {1{`RANDOM}};
  r_907 = _RAND_907[0:0];
  _RAND_908 = {1{`RANDOM}};
  r_908 = _RAND_908[0:0];
  _RAND_909 = {1{`RANDOM}};
  r_909 = _RAND_909[0:0];
  _RAND_910 = {1{`RANDOM}};
  r_910 = _RAND_910[0:0];
  _RAND_911 = {1{`RANDOM}};
  r_911 = _RAND_911[0:0];
  _RAND_912 = {1{`RANDOM}};
  r_912 = _RAND_912[0:0];
  _RAND_913 = {1{`RANDOM}};
  r_913 = _RAND_913[0:0];
  _RAND_914 = {1{`RANDOM}};
  r_914 = _RAND_914[0:0];
  _RAND_915 = {1{`RANDOM}};
  r_915 = _RAND_915[0:0];
  _RAND_916 = {1{`RANDOM}};
  r_916 = _RAND_916[0:0];
  _RAND_917 = {1{`RANDOM}};
  r_917 = _RAND_917[0:0];
  _RAND_918 = {1{`RANDOM}};
  r_918 = _RAND_918[0:0];
  _RAND_919 = {1{`RANDOM}};
  r_919 = _RAND_919[0:0];
  _RAND_920 = {1{`RANDOM}};
  r_920 = _RAND_920[0:0];
  _RAND_921 = {1{`RANDOM}};
  r_921 = _RAND_921[0:0];
  _RAND_922 = {1{`RANDOM}};
  r_922 = _RAND_922[0:0];
  _RAND_923 = {1{`RANDOM}};
  r_923 = _RAND_923[0:0];
  _RAND_924 = {1{`RANDOM}};
  r_924 = _RAND_924[0:0];
  _RAND_925 = {1{`RANDOM}};
  r_925 = _RAND_925[0:0];
  _RAND_926 = {1{`RANDOM}};
  r_926 = _RAND_926[0:0];
  _RAND_927 = {1{`RANDOM}};
  r_927 = _RAND_927[0:0];
  _RAND_928 = {1{`RANDOM}};
  r_928 = _RAND_928[0:0];
  _RAND_929 = {1{`RANDOM}};
  r_929 = _RAND_929[0:0];
  _RAND_930 = {1{`RANDOM}};
  r_930 = _RAND_930[0:0];
  _RAND_931 = {1{`RANDOM}};
  r_931 = _RAND_931[0:0];
  _RAND_932 = {1{`RANDOM}};
  r_932 = _RAND_932[0:0];
  _RAND_933 = {1{`RANDOM}};
  r_933 = _RAND_933[0:0];
  _RAND_934 = {1{`RANDOM}};
  r_934 = _RAND_934[0:0];
  _RAND_935 = {1{`RANDOM}};
  r_935 = _RAND_935[0:0];
  _RAND_936 = {1{`RANDOM}};
  r_936 = _RAND_936[0:0];
  _RAND_937 = {1{`RANDOM}};
  r_937 = _RAND_937[0:0];
  _RAND_938 = {1{`RANDOM}};
  r_938 = _RAND_938[0:0];
  _RAND_939 = {1{`RANDOM}};
  r_939 = _RAND_939[0:0];
  _RAND_940 = {1{`RANDOM}};
  r_940 = _RAND_940[0:0];
  _RAND_941 = {1{`RANDOM}};
  r_941 = _RAND_941[0:0];
  _RAND_942 = {1{`RANDOM}};
  r_942 = _RAND_942[0:0];
  _RAND_943 = {1{`RANDOM}};
  r_943 = _RAND_943[0:0];
  _RAND_944 = {1{`RANDOM}};
  r_944 = _RAND_944[0:0];
  _RAND_945 = {1{`RANDOM}};
  r_945 = _RAND_945[0:0];
  _RAND_946 = {1{`RANDOM}};
  r_946 = _RAND_946[0:0];
  _RAND_947 = {1{`RANDOM}};
  r_947 = _RAND_947[0:0];
  _RAND_948 = {1{`RANDOM}};
  r_948 = _RAND_948[0:0];
  _RAND_949 = {1{`RANDOM}};
  r_949 = _RAND_949[0:0];
  _RAND_950 = {1{`RANDOM}};
  r_950 = _RAND_950[0:0];
  _RAND_951 = {1{`RANDOM}};
  r_951 = _RAND_951[0:0];
  _RAND_952 = {1{`RANDOM}};
  r_952 = _RAND_952[0:0];
  _RAND_953 = {1{`RANDOM}};
  r_953 = _RAND_953[0:0];
  _RAND_954 = {1{`RANDOM}};
  r_954 = _RAND_954[0:0];
  _RAND_955 = {1{`RANDOM}};
  r_955 = _RAND_955[0:0];
  _RAND_956 = {1{`RANDOM}};
  r_956 = _RAND_956[0:0];
  _RAND_957 = {1{`RANDOM}};
  r_957 = _RAND_957[0:0];
  _RAND_958 = {1{`RANDOM}};
  r_958 = _RAND_958[0:0];
  _RAND_959 = {1{`RANDOM}};
  r_959 = _RAND_959[0:0];
  _RAND_960 = {1{`RANDOM}};
  r_960 = _RAND_960[0:0];
  _RAND_961 = {1{`RANDOM}};
  r_961 = _RAND_961[0:0];
  _RAND_962 = {1{`RANDOM}};
  r_962 = _RAND_962[0:0];
  _RAND_963 = {1{`RANDOM}};
  r_963 = _RAND_963[0:0];
  _RAND_964 = {1{`RANDOM}};
  r_964 = _RAND_964[0:0];
  _RAND_965 = {1{`RANDOM}};
  r_965 = _RAND_965[0:0];
  _RAND_966 = {1{`RANDOM}};
  r_966 = _RAND_966[0:0];
  _RAND_967 = {1{`RANDOM}};
  r_967 = _RAND_967[0:0];
  _RAND_968 = {1{`RANDOM}};
  r_968 = _RAND_968[0:0];
  _RAND_969 = {1{`RANDOM}};
  r_969 = _RAND_969[0:0];
  _RAND_970 = {1{`RANDOM}};
  r_970 = _RAND_970[0:0];
  _RAND_971 = {1{`RANDOM}};
  r_971 = _RAND_971[0:0];
  _RAND_972 = {1{`RANDOM}};
  r_972 = _RAND_972[0:0];
  _RAND_973 = {1{`RANDOM}};
  r_973 = _RAND_973[0:0];
  _RAND_974 = {1{`RANDOM}};
  r_974 = _RAND_974[0:0];
  _RAND_975 = {1{`RANDOM}};
  r_975 = _RAND_975[0:0];
  _RAND_976 = {1{`RANDOM}};
  r_976 = _RAND_976[0:0];
  _RAND_977 = {1{`RANDOM}};
  r_977 = _RAND_977[0:0];
  _RAND_978 = {1{`RANDOM}};
  r_978 = _RAND_978[0:0];
  _RAND_979 = {1{`RANDOM}};
  r_979 = _RAND_979[0:0];
  _RAND_980 = {1{`RANDOM}};
  r_980 = _RAND_980[0:0];
  _RAND_981 = {1{`RANDOM}};
  r_981 = _RAND_981[0:0];
  _RAND_982 = {1{`RANDOM}};
  r_982 = _RAND_982[0:0];
  _RAND_983 = {1{`RANDOM}};
  r_983 = _RAND_983[0:0];
  _RAND_984 = {1{`RANDOM}};
  r_984 = _RAND_984[0:0];
  _RAND_985 = {1{`RANDOM}};
  r_985 = _RAND_985[0:0];
  _RAND_986 = {1{`RANDOM}};
  r_986 = _RAND_986[0:0];
  _RAND_987 = {1{`RANDOM}};
  r_987 = _RAND_987[0:0];
  _RAND_988 = {1{`RANDOM}};
  r_988 = _RAND_988[0:0];
  _RAND_989 = {1{`RANDOM}};
  r_989 = _RAND_989[0:0];
  _RAND_990 = {1{`RANDOM}};
  r_990 = _RAND_990[0:0];
  _RAND_991 = {1{`RANDOM}};
  r_991 = _RAND_991[0:0];
  _RAND_992 = {1{`RANDOM}};
  r_992 = _RAND_992[0:0];
  _RAND_993 = {1{`RANDOM}};
  r_993 = _RAND_993[0:0];
  _RAND_994 = {1{`RANDOM}};
  r_994 = _RAND_994[0:0];
  _RAND_995 = {1{`RANDOM}};
  r_995 = _RAND_995[0:0];
  _RAND_996 = {1{`RANDOM}};
  r_996 = _RAND_996[0:0];
  _RAND_997 = {1{`RANDOM}};
  r_997 = _RAND_997[0:0];
  _RAND_998 = {1{`RANDOM}};
  r_998 = _RAND_998[0:0];
  _RAND_999 = {1{`RANDOM}};
  r_999 = _RAND_999[0:0];
  _RAND_1000 = {1{`RANDOM}};
  r_1000 = _RAND_1000[0:0];
  _RAND_1001 = {1{`RANDOM}};
  r_1001 = _RAND_1001[0:0];
  _RAND_1002 = {1{`RANDOM}};
  r_1002 = _RAND_1002[0:0];
  _RAND_1003 = {1{`RANDOM}};
  r_1003 = _RAND_1003[0:0];
  _RAND_1004 = {1{`RANDOM}};
  r_1004 = _RAND_1004[0:0];
  _RAND_1005 = {1{`RANDOM}};
  r_1005 = _RAND_1005[0:0];
  _RAND_1006 = {1{`RANDOM}};
  r_1006 = _RAND_1006[0:0];
  _RAND_1007 = {1{`RANDOM}};
  r_1007 = _RAND_1007[0:0];
  _RAND_1008 = {1{`RANDOM}};
  r_1008 = _RAND_1008[0:0];
  _RAND_1009 = {1{`RANDOM}};
  r_1009 = _RAND_1009[0:0];
  _RAND_1010 = {1{`RANDOM}};
  r_1010 = _RAND_1010[0:0];
  _RAND_1011 = {1{`RANDOM}};
  r_1011 = _RAND_1011[0:0];
  _RAND_1012 = {1{`RANDOM}};
  r_1012 = _RAND_1012[0:0];
  _RAND_1013 = {1{`RANDOM}};
  r_1013 = _RAND_1013[0:0];
  _RAND_1014 = {1{`RANDOM}};
  r_1014 = _RAND_1014[0:0];
  _RAND_1015 = {1{`RANDOM}};
  r_1015 = _RAND_1015[0:0];
  _RAND_1016 = {1{`RANDOM}};
  r_1016 = _RAND_1016[0:0];
  _RAND_1017 = {1{`RANDOM}};
  r_1017 = _RAND_1017[0:0];
  _RAND_1018 = {1{`RANDOM}};
  r_1018 = _RAND_1018[0:0];
  _RAND_1019 = {1{`RANDOM}};
  r_1019 = _RAND_1019[0:0];
  _RAND_1020 = {1{`RANDOM}};
  r_1020 = _RAND_1020[0:0];
  _RAND_1021 = {1{`RANDOM}};
  r_1021 = _RAND_1021[0:0];
  _RAND_1022 = {1{`RANDOM}};
  r_1022 = _RAND_1022[0:0];
  _RAND_1023 = {1{`RANDOM}};
  r_1023 = _RAND_1023[0:0];
  _RAND_1024 = {1{`RANDOM}};
  r_1024 = _RAND_1024[0:0];
  _RAND_1025 = {1{`RANDOM}};
  r_1025 = _RAND_1025[0:0];
  _RAND_1026 = {1{`RANDOM}};
  r_1026 = _RAND_1026[0:0];
  _RAND_1027 = {1{`RANDOM}};
  r_1027 = _RAND_1027[0:0];
  _RAND_1028 = {1{`RANDOM}};
  r_1028 = _RAND_1028[0:0];
  _RAND_1029 = {1{`RANDOM}};
  r_1029 = _RAND_1029[0:0];
  _RAND_1030 = {1{`RANDOM}};
  r_1030 = _RAND_1030[0:0];
  _RAND_1031 = {1{`RANDOM}};
  r_1031 = _RAND_1031[0:0];
  _RAND_1032 = {1{`RANDOM}};
  r_1032 = _RAND_1032[0:0];
  _RAND_1033 = {1{`RANDOM}};
  r_1033 = _RAND_1033[0:0];
  _RAND_1034 = {1{`RANDOM}};
  r_1034 = _RAND_1034[0:0];
  _RAND_1035 = {1{`RANDOM}};
  r_1035 = _RAND_1035[0:0];
  _RAND_1036 = {1{`RANDOM}};
  r_1036 = _RAND_1036[0:0];
  _RAND_1037 = {1{`RANDOM}};
  r_1037 = _RAND_1037[0:0];
  _RAND_1038 = {1{`RANDOM}};
  r_1038 = _RAND_1038[0:0];
  _RAND_1039 = {1{`RANDOM}};
  r_1039 = _RAND_1039[0:0];
  _RAND_1040 = {1{`RANDOM}};
  r_1040 = _RAND_1040[0:0];
  _RAND_1041 = {1{`RANDOM}};
  r_1041 = _RAND_1041[0:0];
  _RAND_1042 = {1{`RANDOM}};
  r_1042 = _RAND_1042[0:0];
  _RAND_1043 = {1{`RANDOM}};
  r_1043 = _RAND_1043[0:0];
  _RAND_1044 = {1{`RANDOM}};
  r_1044 = _RAND_1044[0:0];
  _RAND_1045 = {1{`RANDOM}};
  r_1045 = _RAND_1045[0:0];
  _RAND_1046 = {1{`RANDOM}};
  r_1046 = _RAND_1046[0:0];
  _RAND_1047 = {1{`RANDOM}};
  r_1047 = _RAND_1047[0:0];
  _RAND_1048 = {1{`RANDOM}};
  r_1048 = _RAND_1048[0:0];
  _RAND_1049 = {1{`RANDOM}};
  r_1049 = _RAND_1049[0:0];
  _RAND_1050 = {1{`RANDOM}};
  r_1050 = _RAND_1050[0:0];
  _RAND_1051 = {1{`RANDOM}};
  r_1051 = _RAND_1051[0:0];
  _RAND_1052 = {1{`RANDOM}};
  r_1052 = _RAND_1052[0:0];
  _RAND_1053 = {1{`RANDOM}};
  r_1053 = _RAND_1053[0:0];
  _RAND_1054 = {1{`RANDOM}};
  r_1054 = _RAND_1054[0:0];
  _RAND_1055 = {1{`RANDOM}};
  r_1055 = _RAND_1055[0:0];
  _RAND_1056 = {1{`RANDOM}};
  r_1056 = _RAND_1056[0:0];
  _RAND_1057 = {1{`RANDOM}};
  r_1057 = _RAND_1057[0:0];
  _RAND_1058 = {1{`RANDOM}};
  r_1058 = _RAND_1058[0:0];
  _RAND_1059 = {1{`RANDOM}};
  r_1059 = _RAND_1059[0:0];
  _RAND_1060 = {1{`RANDOM}};
  r_1060 = _RAND_1060[0:0];
  _RAND_1061 = {1{`RANDOM}};
  r_1061 = _RAND_1061[0:0];
  _RAND_1062 = {1{`RANDOM}};
  r_1062 = _RAND_1062[0:0];
  _RAND_1063 = {1{`RANDOM}};
  r_1063 = _RAND_1063[0:0];
  _RAND_1064 = {1{`RANDOM}};
  r_1064 = _RAND_1064[0:0];
  _RAND_1065 = {1{`RANDOM}};
  r_1065 = _RAND_1065[0:0];
  _RAND_1066 = {1{`RANDOM}};
  r_1066 = _RAND_1066[0:0];
  _RAND_1067 = {1{`RANDOM}};
  r_1067 = _RAND_1067[0:0];
  _RAND_1068 = {1{`RANDOM}};
  r_1068 = _RAND_1068[0:0];
  _RAND_1069 = {1{`RANDOM}};
  r_1069 = _RAND_1069[0:0];
  _RAND_1070 = {1{`RANDOM}};
  r_1070 = _RAND_1070[0:0];
  _RAND_1071 = {1{`RANDOM}};
  r_1071 = _RAND_1071[0:0];
  _RAND_1072 = {1{`RANDOM}};
  r_1072 = _RAND_1072[0:0];
  _RAND_1073 = {1{`RANDOM}};
  r_1073 = _RAND_1073[0:0];
  _RAND_1074 = {1{`RANDOM}};
  r_1074 = _RAND_1074[0:0];
  _RAND_1075 = {1{`RANDOM}};
  r_1075 = _RAND_1075[0:0];
  _RAND_1076 = {1{`RANDOM}};
  r_1076 = _RAND_1076[0:0];
  _RAND_1077 = {1{`RANDOM}};
  r_1077 = _RAND_1077[0:0];
  _RAND_1078 = {1{`RANDOM}};
  r_1078 = _RAND_1078[0:0];
  _RAND_1079 = {1{`RANDOM}};
  r_1079 = _RAND_1079[0:0];
  _RAND_1080 = {1{`RANDOM}};
  r_1080 = _RAND_1080[0:0];
  _RAND_1081 = {1{`RANDOM}};
  r_1081 = _RAND_1081[0:0];
  _RAND_1082 = {1{`RANDOM}};
  r_1082 = _RAND_1082[0:0];
  _RAND_1083 = {1{`RANDOM}};
  r_1083 = _RAND_1083[0:0];
  _RAND_1084 = {1{`RANDOM}};
  r_1084 = _RAND_1084[0:0];
  _RAND_1085 = {1{`RANDOM}};
  r_1085 = _RAND_1085[0:0];
  _RAND_1086 = {1{`RANDOM}};
  r_1086 = _RAND_1086[0:0];
  _RAND_1087 = {1{`RANDOM}};
  r_1087 = _RAND_1087[0:0];
  _RAND_1088 = {1{`RANDOM}};
  r_1088 = _RAND_1088[0:0];
  _RAND_1089 = {1{`RANDOM}};
  r_1089 = _RAND_1089[0:0];
  _RAND_1090 = {1{`RANDOM}};
  r_1090 = _RAND_1090[0:0];
  _RAND_1091 = {1{`RANDOM}};
  r_1091 = _RAND_1091[0:0];
  _RAND_1092 = {1{`RANDOM}};
  r_1092 = _RAND_1092[0:0];
  _RAND_1093 = {1{`RANDOM}};
  r_1093 = _RAND_1093[0:0];
  _RAND_1094 = {1{`RANDOM}};
  r_1094 = _RAND_1094[0:0];
  _RAND_1095 = {1{`RANDOM}};
  r_1095 = _RAND_1095[0:0];
  _RAND_1096 = {1{`RANDOM}};
  r_1096 = _RAND_1096[0:0];
  _RAND_1097 = {1{`RANDOM}};
  r_1097 = _RAND_1097[0:0];
  _RAND_1098 = {1{`RANDOM}};
  r_1098 = _RAND_1098[0:0];
  _RAND_1099 = {1{`RANDOM}};
  r_1099 = _RAND_1099[0:0];
  _RAND_1100 = {1{`RANDOM}};
  r_1100 = _RAND_1100[0:0];
  _RAND_1101 = {1{`RANDOM}};
  r_1101 = _RAND_1101[0:0];
  _RAND_1102 = {1{`RANDOM}};
  r_1102 = _RAND_1102[0:0];
  _RAND_1103 = {1{`RANDOM}};
  r_1103 = _RAND_1103[0:0];
  _RAND_1104 = {1{`RANDOM}};
  r_1104 = _RAND_1104[0:0];
  _RAND_1105 = {1{`RANDOM}};
  r_1105 = _RAND_1105[0:0];
  _RAND_1106 = {1{`RANDOM}};
  r_1106 = _RAND_1106[0:0];
  _RAND_1107 = {1{`RANDOM}};
  r_1107 = _RAND_1107[0:0];
  _RAND_1108 = {1{`RANDOM}};
  r_1108 = _RAND_1108[0:0];
  _RAND_1109 = {1{`RANDOM}};
  r_1109 = _RAND_1109[0:0];
  _RAND_1110 = {1{`RANDOM}};
  r_1110 = _RAND_1110[0:0];
  _RAND_1111 = {1{`RANDOM}};
  r_1111 = _RAND_1111[0:0];
  _RAND_1112 = {1{`RANDOM}};
  r_1112 = _RAND_1112[0:0];
  _RAND_1113 = {1{`RANDOM}};
  r_1113 = _RAND_1113[0:0];
  _RAND_1114 = {1{`RANDOM}};
  r_1114 = _RAND_1114[0:0];
  _RAND_1115 = {1{`RANDOM}};
  r_1115 = _RAND_1115[0:0];
  _RAND_1116 = {1{`RANDOM}};
  r_1116 = _RAND_1116[0:0];
  _RAND_1117 = {1{`RANDOM}};
  r_1117 = _RAND_1117[0:0];
  _RAND_1118 = {1{`RANDOM}};
  r_1118 = _RAND_1118[0:0];
  _RAND_1119 = {1{`RANDOM}};
  r_1119 = _RAND_1119[0:0];
  _RAND_1120 = {1{`RANDOM}};
  r_1120 = _RAND_1120[0:0];
  _RAND_1121 = {1{`RANDOM}};
  r_1121 = _RAND_1121[0:0];
  _RAND_1122 = {1{`RANDOM}};
  r_1122 = _RAND_1122[0:0];
  _RAND_1123 = {1{`RANDOM}};
  r_1123 = _RAND_1123[0:0];
  _RAND_1124 = {1{`RANDOM}};
  r_1124 = _RAND_1124[0:0];
  _RAND_1125 = {1{`RANDOM}};
  r_1125 = _RAND_1125[0:0];
  _RAND_1126 = {1{`RANDOM}};
  r_1126 = _RAND_1126[0:0];
  _RAND_1127 = {1{`RANDOM}};
  r_1127 = _RAND_1127[0:0];
  _RAND_1128 = {1{`RANDOM}};
  r_1128 = _RAND_1128[0:0];
  _RAND_1129 = {1{`RANDOM}};
  r_1129 = _RAND_1129[0:0];
  _RAND_1130 = {1{`RANDOM}};
  r_1130 = _RAND_1130[0:0];
  _RAND_1131 = {1{`RANDOM}};
  r_1131 = _RAND_1131[0:0];
  _RAND_1132 = {1{`RANDOM}};
  r_1132 = _RAND_1132[0:0];
  _RAND_1133 = {1{`RANDOM}};
  r_1133 = _RAND_1133[0:0];
  _RAND_1134 = {1{`RANDOM}};
  r_1134 = _RAND_1134[0:0];
  _RAND_1135 = {1{`RANDOM}};
  r_1135 = _RAND_1135[0:0];
  _RAND_1136 = {1{`RANDOM}};
  r_1136 = _RAND_1136[0:0];
  _RAND_1137 = {1{`RANDOM}};
  r_1137 = _RAND_1137[0:0];
  _RAND_1138 = {1{`RANDOM}};
  r_1138 = _RAND_1138[0:0];
  _RAND_1139 = {1{`RANDOM}};
  r_1139 = _RAND_1139[0:0];
  _RAND_1140 = {1{`RANDOM}};
  r_1140 = _RAND_1140[0:0];
  _RAND_1141 = {1{`RANDOM}};
  r_1141 = _RAND_1141[0:0];
  _RAND_1142 = {1{`RANDOM}};
  r_1142 = _RAND_1142[0:0];
  _RAND_1143 = {1{`RANDOM}};
  r_1143 = _RAND_1143[0:0];
  _RAND_1144 = {1{`RANDOM}};
  r_1144 = _RAND_1144[0:0];
  _RAND_1145 = {1{`RANDOM}};
  r_1145 = _RAND_1145[0:0];
  _RAND_1146 = {1{`RANDOM}};
  r_1146 = _RAND_1146[0:0];
  _RAND_1147 = {1{`RANDOM}};
  r_1147 = _RAND_1147[0:0];
  _RAND_1148 = {1{`RANDOM}};
  r_1148 = _RAND_1148[0:0];
  _RAND_1149 = {1{`RANDOM}};
  r_1149 = _RAND_1149[0:0];
  _RAND_1150 = {1{`RANDOM}};
  r_1150 = _RAND_1150[0:0];
  _RAND_1151 = {1{`RANDOM}};
  r_1151 = _RAND_1151[0:0];
  _RAND_1152 = {1{`RANDOM}};
  r_1152 = _RAND_1152[0:0];
  _RAND_1153 = {1{`RANDOM}};
  r_1153 = _RAND_1153[0:0];
  _RAND_1154 = {1{`RANDOM}};
  r_1154 = _RAND_1154[0:0];
  _RAND_1155 = {1{`RANDOM}};
  r_1155 = _RAND_1155[0:0];
  _RAND_1156 = {1{`RANDOM}};
  r_1156 = _RAND_1156[0:0];
  _RAND_1157 = {1{`RANDOM}};
  r_1157 = _RAND_1157[0:0];
  _RAND_1158 = {1{`RANDOM}};
  r_1158 = _RAND_1158[0:0];
  _RAND_1159 = {1{`RANDOM}};
  r_1159 = _RAND_1159[0:0];
  _RAND_1160 = {1{`RANDOM}};
  r_1160 = _RAND_1160[0:0];
  _RAND_1161 = {1{`RANDOM}};
  r_1161 = _RAND_1161[0:0];
  _RAND_1162 = {1{`RANDOM}};
  r_1162 = _RAND_1162[0:0];
  _RAND_1163 = {1{`RANDOM}};
  r_1163 = _RAND_1163[0:0];
  _RAND_1164 = {1{`RANDOM}};
  r_1164 = _RAND_1164[0:0];
  _RAND_1165 = {1{`RANDOM}};
  r_1165 = _RAND_1165[0:0];
  _RAND_1166 = {1{`RANDOM}};
  r_1166 = _RAND_1166[0:0];
  _RAND_1167 = {1{`RANDOM}};
  r_1167 = _RAND_1167[0:0];
  _RAND_1168 = {1{`RANDOM}};
  r_1168 = _RAND_1168[0:0];
  _RAND_1169 = {1{`RANDOM}};
  r_1169 = _RAND_1169[0:0];
  _RAND_1170 = {1{`RANDOM}};
  r_1170 = _RAND_1170[0:0];
  _RAND_1171 = {1{`RANDOM}};
  r_1171 = _RAND_1171[0:0];
  _RAND_1172 = {1{`RANDOM}};
  r_1172 = _RAND_1172[0:0];
  _RAND_1173 = {1{`RANDOM}};
  r_1173 = _RAND_1173[0:0];
  _RAND_1174 = {1{`RANDOM}};
  r_1174 = _RAND_1174[0:0];
  _RAND_1175 = {1{`RANDOM}};
  r_1175 = _RAND_1175[0:0];
  _RAND_1176 = {1{`RANDOM}};
  r_1176 = _RAND_1176[0:0];
  _RAND_1177 = {1{`RANDOM}};
  r_1177 = _RAND_1177[0:0];
  _RAND_1178 = {1{`RANDOM}};
  r_1178 = _RAND_1178[0:0];
  _RAND_1179 = {1{`RANDOM}};
  r_1179 = _RAND_1179[0:0];
  _RAND_1180 = {1{`RANDOM}};
  r_1180 = _RAND_1180[0:0];
  _RAND_1181 = {1{`RANDOM}};
  r_1181 = _RAND_1181[0:0];
  _RAND_1182 = {1{`RANDOM}};
  r_1182 = _RAND_1182[0:0];
  _RAND_1183 = {1{`RANDOM}};
  r_1183 = _RAND_1183[0:0];
  _RAND_1184 = {1{`RANDOM}};
  r_1184 = _RAND_1184[0:0];
  _RAND_1185 = {1{`RANDOM}};
  r_1185 = _RAND_1185[0:0];
  _RAND_1186 = {1{`RANDOM}};
  r_1186 = _RAND_1186[0:0];
  _RAND_1187 = {1{`RANDOM}};
  r_1187 = _RAND_1187[0:0];
  _RAND_1188 = {1{`RANDOM}};
  r_1188 = _RAND_1188[0:0];
  _RAND_1189 = {1{`RANDOM}};
  r_1189 = _RAND_1189[0:0];
  _RAND_1190 = {1{`RANDOM}};
  r_1190 = _RAND_1190[0:0];
  _RAND_1191 = {1{`RANDOM}};
  r_1191 = _RAND_1191[0:0];
  _RAND_1192 = {1{`RANDOM}};
  r_1192 = _RAND_1192[0:0];
  _RAND_1193 = {1{`RANDOM}};
  r_1193 = _RAND_1193[0:0];
  _RAND_1194 = {1{`RANDOM}};
  r_1194 = _RAND_1194[0:0];
  _RAND_1195 = {1{`RANDOM}};
  r_1195 = _RAND_1195[0:0];
  _RAND_1196 = {1{`RANDOM}};
  r_1196 = _RAND_1196[0:0];
  _RAND_1197 = {1{`RANDOM}};
  r_1197 = _RAND_1197[0:0];
  _RAND_1198 = {1{`RANDOM}};
  r_1198 = _RAND_1198[0:0];
  _RAND_1199 = {1{`RANDOM}};
  r_1199 = _RAND_1199[0:0];
  _RAND_1200 = {1{`RANDOM}};
  r_1200 = _RAND_1200[0:0];
  _RAND_1201 = {1{`RANDOM}};
  r_1201 = _RAND_1201[0:0];
  _RAND_1202 = {1{`RANDOM}};
  r_1202 = _RAND_1202[0:0];
  _RAND_1203 = {1{`RANDOM}};
  r_1203 = _RAND_1203[0:0];
  _RAND_1204 = {1{`RANDOM}};
  r_1204 = _RAND_1204[0:0];
  _RAND_1205 = {1{`RANDOM}};
  r_1205 = _RAND_1205[0:0];
  _RAND_1206 = {1{`RANDOM}};
  r_1206 = _RAND_1206[0:0];
  _RAND_1207 = {1{`RANDOM}};
  r_1207 = _RAND_1207[0:0];
  _RAND_1208 = {1{`RANDOM}};
  r_1208 = _RAND_1208[0:0];
  _RAND_1209 = {1{`RANDOM}};
  r_1209 = _RAND_1209[0:0];
  _RAND_1210 = {1{`RANDOM}};
  r_1210 = _RAND_1210[0:0];
  _RAND_1211 = {1{`RANDOM}};
  r_1211 = _RAND_1211[0:0];
  _RAND_1212 = {1{`RANDOM}};
  r_1212 = _RAND_1212[0:0];
  _RAND_1213 = {1{`RANDOM}};
  r_1213 = _RAND_1213[0:0];
  _RAND_1214 = {1{`RANDOM}};
  r_1214 = _RAND_1214[0:0];
  _RAND_1215 = {1{`RANDOM}};
  r_1215 = _RAND_1215[0:0];
  _RAND_1216 = {1{`RANDOM}};
  r_1216 = _RAND_1216[0:0];
  _RAND_1217 = {1{`RANDOM}};
  r_1217 = _RAND_1217[0:0];
  _RAND_1218 = {1{`RANDOM}};
  r_1218 = _RAND_1218[0:0];
  _RAND_1219 = {1{`RANDOM}};
  r_1219 = _RAND_1219[0:0];
  _RAND_1220 = {1{`RANDOM}};
  r_1220 = _RAND_1220[0:0];
  _RAND_1221 = {1{`RANDOM}};
  r_1221 = _RAND_1221[0:0];
  _RAND_1222 = {1{`RANDOM}};
  r_1222 = _RAND_1222[0:0];
  _RAND_1223 = {1{`RANDOM}};
  r_1223 = _RAND_1223[0:0];
  _RAND_1224 = {1{`RANDOM}};
  r_1224 = _RAND_1224[0:0];
  _RAND_1225 = {1{`RANDOM}};
  r_1225 = _RAND_1225[0:0];
  _RAND_1226 = {1{`RANDOM}};
  r_1226 = _RAND_1226[0:0];
  _RAND_1227 = {1{`RANDOM}};
  r_1227 = _RAND_1227[0:0];
  _RAND_1228 = {1{`RANDOM}};
  r_1228 = _RAND_1228[0:0];
  _RAND_1229 = {1{`RANDOM}};
  r_1229 = _RAND_1229[0:0];
  _RAND_1230 = {1{`RANDOM}};
  r_1230 = _RAND_1230[0:0];
  _RAND_1231 = {1{`RANDOM}};
  r_1231 = _RAND_1231[0:0];
  _RAND_1232 = {1{`RANDOM}};
  r_1232 = _RAND_1232[0:0];
  _RAND_1233 = {1{`RANDOM}};
  r_1233 = _RAND_1233[0:0];
  _RAND_1234 = {1{`RANDOM}};
  r_1234 = _RAND_1234[0:0];
  _RAND_1235 = {1{`RANDOM}};
  r_1235 = _RAND_1235[0:0];
  _RAND_1236 = {1{`RANDOM}};
  r_1236 = _RAND_1236[0:0];
  _RAND_1237 = {1{`RANDOM}};
  r_1237 = _RAND_1237[0:0];
  _RAND_1238 = {1{`RANDOM}};
  r_1238 = _RAND_1238[0:0];
  _RAND_1239 = {1{`RANDOM}};
  r_1239 = _RAND_1239[0:0];
  _RAND_1240 = {1{`RANDOM}};
  r_1240 = _RAND_1240[0:0];
  _RAND_1241 = {1{`RANDOM}};
  r_1241 = _RAND_1241[0:0];
  _RAND_1242 = {1{`RANDOM}};
  r_1242 = _RAND_1242[0:0];
  _RAND_1243 = {1{`RANDOM}};
  r_1243 = _RAND_1243[0:0];
  _RAND_1244 = {1{`RANDOM}};
  r_1244 = _RAND_1244[0:0];
  _RAND_1245 = {1{`RANDOM}};
  r_1245 = _RAND_1245[0:0];
  _RAND_1246 = {1{`RANDOM}};
  r_1246 = _RAND_1246[0:0];
  _RAND_1247 = {1{`RANDOM}};
  r_1247 = _RAND_1247[0:0];
  _RAND_1248 = {1{`RANDOM}};
  r_1248 = _RAND_1248[0:0];
  _RAND_1249 = {1{`RANDOM}};
  r_1249 = _RAND_1249[0:0];
  _RAND_1250 = {1{`RANDOM}};
  r_1250 = _RAND_1250[0:0];
  _RAND_1251 = {1{`RANDOM}};
  r_1251 = _RAND_1251[0:0];
  _RAND_1252 = {1{`RANDOM}};
  r_1252 = _RAND_1252[0:0];
  _RAND_1253 = {1{`RANDOM}};
  r_1253 = _RAND_1253[0:0];
  _RAND_1254 = {1{`RANDOM}};
  r_1254 = _RAND_1254[0:0];
  _RAND_1255 = {1{`RANDOM}};
  r_1255 = _RAND_1255[0:0];
  _RAND_1256 = {1{`RANDOM}};
  r_1256 = _RAND_1256[0:0];
  _RAND_1257 = {1{`RANDOM}};
  r_1257 = _RAND_1257[0:0];
  _RAND_1258 = {1{`RANDOM}};
  r_1258 = _RAND_1258[0:0];
  _RAND_1259 = {1{`RANDOM}};
  r_1259 = _RAND_1259[0:0];
  _RAND_1260 = {1{`RANDOM}};
  r_1260 = _RAND_1260[0:0];
  _RAND_1261 = {1{`RANDOM}};
  r_1261 = _RAND_1261[0:0];
  _RAND_1262 = {1{`RANDOM}};
  r_1262 = _RAND_1262[0:0];
  _RAND_1263 = {1{`RANDOM}};
  r_1263 = _RAND_1263[0:0];
  _RAND_1264 = {1{`RANDOM}};
  r_1264 = _RAND_1264[0:0];
  _RAND_1265 = {1{`RANDOM}};
  r_1265 = _RAND_1265[0:0];
  _RAND_1266 = {1{`RANDOM}};
  r_1266 = _RAND_1266[0:0];
  _RAND_1267 = {1{`RANDOM}};
  r_1267 = _RAND_1267[0:0];
  _RAND_1268 = {1{`RANDOM}};
  r_1268 = _RAND_1268[0:0];
  _RAND_1269 = {1{`RANDOM}};
  r_1269 = _RAND_1269[0:0];
  _RAND_1270 = {1{`RANDOM}};
  r_1270 = _RAND_1270[0:0];
  _RAND_1271 = {1{`RANDOM}};
  r_1271 = _RAND_1271[0:0];
  _RAND_1272 = {1{`RANDOM}};
  r_1272 = _RAND_1272[0:0];
  _RAND_1273 = {1{`RANDOM}};
  r_1273 = _RAND_1273[0:0];
  _RAND_1274 = {1{`RANDOM}};
  r_1274 = _RAND_1274[0:0];
  _RAND_1275 = {1{`RANDOM}};
  r_1275 = _RAND_1275[0:0];
  _RAND_1276 = {1{`RANDOM}};
  r_1276 = _RAND_1276[0:0];
  _RAND_1277 = {1{`RANDOM}};
  r_1277 = _RAND_1277[0:0];
  _RAND_1278 = {1{`RANDOM}};
  r_1278 = _RAND_1278[0:0];
  _RAND_1279 = {1{`RANDOM}};
  r_1279 = _RAND_1279[0:0];
  _RAND_1280 = {1{`RANDOM}};
  r_1280 = _RAND_1280[0:0];
  _RAND_1281 = {1{`RANDOM}};
  r_1281 = _RAND_1281[0:0];
  _RAND_1282 = {1{`RANDOM}};
  r_1282 = _RAND_1282[0:0];
  _RAND_1283 = {1{`RANDOM}};
  r_1283 = _RAND_1283[0:0];
  _RAND_1284 = {1{`RANDOM}};
  r_1284 = _RAND_1284[0:0];
  _RAND_1285 = {1{`RANDOM}};
  r_1286 = _RAND_1285[0:0];
  _RAND_1286 = {1{`RANDOM}};
  r_1287 = _RAND_1286[0:0];
  _RAND_1287 = {1{`RANDOM}};
  r_1288 = _RAND_1287[0:0];
  _RAND_1288 = {1{`RANDOM}};
  r_1289 = _RAND_1288[0:0];
  _RAND_1289 = {1{`RANDOM}};
  r_1290 = _RAND_1289[0:0];
  _RAND_1290 = {1{`RANDOM}};
  r_1291 = _RAND_1290[0:0];
  _RAND_1291 = {1{`RANDOM}};
  r_1292 = _RAND_1291[0:0];
  _RAND_1292 = {1{`RANDOM}};
  r_1293 = _RAND_1292[0:0];
  _RAND_1293 = {1{`RANDOM}};
  r_1294 = _RAND_1293[0:0];
  _RAND_1294 = {1{`RANDOM}};
  r_1295 = _RAND_1294[0:0];
  _RAND_1295 = {1{`RANDOM}};
  r_1296 = _RAND_1295[0:0];
  _RAND_1296 = {1{`RANDOM}};
  r_1297 = _RAND_1296[0:0];
  _RAND_1297 = {1{`RANDOM}};
  r_1298 = _RAND_1297[0:0];
  _RAND_1298 = {1{`RANDOM}};
  r_1299 = _RAND_1298[0:0];
  _RAND_1299 = {1{`RANDOM}};
  r_1300 = _RAND_1299[0:0];
  _RAND_1300 = {1{`RANDOM}};
  r_1301 = _RAND_1300[0:0];
  _RAND_1301 = {1{`RANDOM}};
  r_1302 = _RAND_1301[0:0];
  _RAND_1302 = {1{`RANDOM}};
  r_1303 = _RAND_1302[0:0];
  _RAND_1303 = {1{`RANDOM}};
  r_1304 = _RAND_1303[0:0];
  _RAND_1304 = {1{`RANDOM}};
  r_1305 = _RAND_1304[0:0];
  _RAND_1305 = {1{`RANDOM}};
  r_1306 = _RAND_1305[0:0];
  _RAND_1306 = {1{`RANDOM}};
  r_1307 = _RAND_1306[0:0];
  _RAND_1307 = {1{`RANDOM}};
  r_1308 = _RAND_1307[0:0];
  _RAND_1308 = {1{`RANDOM}};
  r_1309 = _RAND_1308[0:0];
  _RAND_1309 = {1{`RANDOM}};
  r_1310 = _RAND_1309[0:0];
  _RAND_1310 = {1{`RANDOM}};
  r_1311 = _RAND_1310[0:0];
  _RAND_1311 = {1{`RANDOM}};
  r_1312 = _RAND_1311[0:0];
  _RAND_1312 = {1{`RANDOM}};
  r_1313 = _RAND_1312[0:0];
  _RAND_1313 = {1{`RANDOM}};
  r_1314 = _RAND_1313[0:0];
  _RAND_1314 = {1{`RANDOM}};
  r_1315 = _RAND_1314[0:0];
  _RAND_1315 = {1{`RANDOM}};
  r_1316 = _RAND_1315[0:0];
  _RAND_1316 = {1{`RANDOM}};
  r_1317 = _RAND_1316[0:0];
  _RAND_1317 = {1{`RANDOM}};
  r_1318 = _RAND_1317[0:0];
  _RAND_1318 = {1{`RANDOM}};
  r_1319 = _RAND_1318[0:0];
  _RAND_1319 = {1{`RANDOM}};
  r_1320 = _RAND_1319[0:0];
  _RAND_1320 = {1{`RANDOM}};
  r_1321 = _RAND_1320[0:0];
  _RAND_1321 = {1{`RANDOM}};
  r_1322 = _RAND_1321[0:0];
  _RAND_1322 = {1{`RANDOM}};
  r_1323 = _RAND_1322[0:0];
  _RAND_1323 = {1{`RANDOM}};
  r_1324 = _RAND_1323[0:0];
  _RAND_1324 = {1{`RANDOM}};
  r_1325 = _RAND_1324[0:0];
  _RAND_1325 = {1{`RANDOM}};
  r_1326 = _RAND_1325[0:0];
  _RAND_1326 = {1{`RANDOM}};
  r_1327 = _RAND_1326[0:0];
  _RAND_1327 = {1{`RANDOM}};
  r_1328 = _RAND_1327[0:0];
  _RAND_1328 = {1{`RANDOM}};
  r_1329 = _RAND_1328[0:0];
  _RAND_1329 = {1{`RANDOM}};
  r_1330 = _RAND_1329[0:0];
  _RAND_1330 = {1{`RANDOM}};
  r_1331 = _RAND_1330[0:0];
  _RAND_1331 = {1{`RANDOM}};
  r_1332 = _RAND_1331[0:0];
  _RAND_1332 = {1{`RANDOM}};
  r_1333 = _RAND_1332[0:0];
  _RAND_1333 = {1{`RANDOM}};
  r_1334 = _RAND_1333[0:0];
  _RAND_1334 = {1{`RANDOM}};
  r_1335 = _RAND_1334[0:0];
  _RAND_1335 = {1{`RANDOM}};
  r_1336 = _RAND_1335[0:0];
  _RAND_1336 = {1{`RANDOM}};
  r_1337 = _RAND_1336[0:0];
  _RAND_1337 = {1{`RANDOM}};
  r_1338 = _RAND_1337[0:0];
  _RAND_1338 = {1{`RANDOM}};
  r_1339 = _RAND_1338[0:0];
  _RAND_1339 = {1{`RANDOM}};
  r_1340 = _RAND_1339[0:0];
  _RAND_1340 = {1{`RANDOM}};
  r_1341 = _RAND_1340[0:0];
  _RAND_1341 = {1{`RANDOM}};
  r_1342 = _RAND_1341[0:0];
  _RAND_1342 = {1{`RANDOM}};
  r_1343 = _RAND_1342[0:0];
  _RAND_1343 = {1{`RANDOM}};
  r_1344 = _RAND_1343[0:0];
  _RAND_1344 = {1{`RANDOM}};
  r_1345 = _RAND_1344[0:0];
  _RAND_1345 = {1{`RANDOM}};
  r_1346 = _RAND_1345[0:0];
  _RAND_1346 = {1{`RANDOM}};
  r_1347 = _RAND_1346[0:0];
  _RAND_1347 = {1{`RANDOM}};
  r_1349 = _RAND_1347[0:0];
  _RAND_1348 = {1{`RANDOM}};
  r_1350 = _RAND_1348[0:0];
  _RAND_1349 = {1{`RANDOM}};
  r_1351 = _RAND_1349[0:0];
  _RAND_1350 = {1{`RANDOM}};
  r_1352 = _RAND_1350[0:0];
  _RAND_1351 = {1{`RANDOM}};
  r_1353 = _RAND_1351[0:0];
  _RAND_1352 = {1{`RANDOM}};
  r_1354 = _RAND_1352[0:0];
  _RAND_1353 = {1{`RANDOM}};
  r_1355 = _RAND_1353[0:0];
  _RAND_1354 = {1{`RANDOM}};
  r_1356 = _RAND_1354[0:0];
  _RAND_1355 = {1{`RANDOM}};
  r_1357 = _RAND_1355[0:0];
  _RAND_1356 = {1{`RANDOM}};
  r_1358 = _RAND_1356[0:0];
  _RAND_1357 = {1{`RANDOM}};
  r_1359 = _RAND_1357[0:0];
  _RAND_1358 = {1{`RANDOM}};
  r_1360 = _RAND_1358[0:0];
  _RAND_1359 = {1{`RANDOM}};
  r_1361 = _RAND_1359[0:0];
  _RAND_1360 = {1{`RANDOM}};
  r_1362 = _RAND_1360[0:0];
  _RAND_1361 = {1{`RANDOM}};
  r_1363 = _RAND_1361[0:0];
  _RAND_1362 = {1{`RANDOM}};
  r_1364 = _RAND_1362[0:0];
  _RAND_1363 = {1{`RANDOM}};
  r_1365 = _RAND_1363[0:0];
  _RAND_1364 = {1{`RANDOM}};
  r_1366 = _RAND_1364[0:0];
  _RAND_1365 = {1{`RANDOM}};
  r_1367 = _RAND_1365[0:0];
  _RAND_1366 = {1{`RANDOM}};
  r_1368 = _RAND_1366[0:0];
  _RAND_1367 = {1{`RANDOM}};
  r_1369 = _RAND_1367[0:0];
  _RAND_1368 = {1{`RANDOM}};
  r_1370 = _RAND_1368[0:0];
  _RAND_1369 = {1{`RANDOM}};
  r_1371 = _RAND_1369[0:0];
  _RAND_1370 = {1{`RANDOM}};
  r_1372 = _RAND_1370[0:0];
  _RAND_1371 = {1{`RANDOM}};
  r_1373 = _RAND_1371[0:0];
  _RAND_1372 = {1{`RANDOM}};
  r_1374 = _RAND_1372[0:0];
  _RAND_1373 = {1{`RANDOM}};
  r_1375 = _RAND_1373[0:0];
  _RAND_1374 = {1{`RANDOM}};
  r_1376 = _RAND_1374[0:0];
  _RAND_1375 = {1{`RANDOM}};
  r_1377 = _RAND_1375[0:0];
  _RAND_1376 = {1{`RANDOM}};
  r_1378 = _RAND_1376[0:0];
  _RAND_1377 = {1{`RANDOM}};
  r_1379 = _RAND_1377[0:0];
  _RAND_1378 = {1{`RANDOM}};
  r_1380 = _RAND_1378[0:0];
  _RAND_1379 = {1{`RANDOM}};
  r_1381 = _RAND_1379[0:0];
  _RAND_1380 = {1{`RANDOM}};
  r_1382 = _RAND_1380[0:0];
  _RAND_1381 = {1{`RANDOM}};
  r_1383 = _RAND_1381[0:0];
  _RAND_1382 = {1{`RANDOM}};
  r_1384 = _RAND_1382[0:0];
  _RAND_1383 = {1{`RANDOM}};
  r_1385 = _RAND_1383[0:0];
  _RAND_1384 = {1{`RANDOM}};
  r_1386 = _RAND_1384[0:0];
  _RAND_1385 = {1{`RANDOM}};
  r_1387 = _RAND_1385[0:0];
  _RAND_1386 = {1{`RANDOM}};
  r_1388 = _RAND_1386[0:0];
  _RAND_1387 = {1{`RANDOM}};
  r_1389 = _RAND_1387[0:0];
  _RAND_1388 = {1{`RANDOM}};
  r_1390 = _RAND_1388[0:0];
  _RAND_1389 = {1{`RANDOM}};
  r_1391 = _RAND_1389[0:0];
  _RAND_1390 = {1{`RANDOM}};
  r_1392 = _RAND_1390[0:0];
  _RAND_1391 = {1{`RANDOM}};
  r_1393 = _RAND_1391[0:0];
  _RAND_1392 = {1{`RANDOM}};
  r_1394 = _RAND_1392[0:0];
  _RAND_1393 = {1{`RANDOM}};
  r_1395 = _RAND_1393[0:0];
  _RAND_1394 = {1{`RANDOM}};
  r_1396 = _RAND_1394[0:0];
  _RAND_1395 = {1{`RANDOM}};
  r_1397 = _RAND_1395[0:0];
  _RAND_1396 = {1{`RANDOM}};
  r_1398 = _RAND_1396[0:0];
  _RAND_1397 = {1{`RANDOM}};
  r_1399 = _RAND_1397[0:0];
  _RAND_1398 = {1{`RANDOM}};
  r_1400 = _RAND_1398[0:0];
  _RAND_1399 = {1{`RANDOM}};
  r_1401 = _RAND_1399[0:0];
  _RAND_1400 = {1{`RANDOM}};
  r_1402 = _RAND_1400[0:0];
  _RAND_1401 = {1{`RANDOM}};
  r_1403 = _RAND_1401[0:0];
  _RAND_1402 = {1{`RANDOM}};
  r_1404 = _RAND_1402[0:0];
  _RAND_1403 = {1{`RANDOM}};
  r_1405 = _RAND_1403[0:0];
  _RAND_1404 = {1{`RANDOM}};
  r_1406 = _RAND_1404[0:0];
  _RAND_1405 = {1{`RANDOM}};
  r_1407 = _RAND_1405[0:0];
  _RAND_1406 = {1{`RANDOM}};
  r_1408 = _RAND_1406[0:0];
  _RAND_1407 = {1{`RANDOM}};
  r_1410 = _RAND_1407[0:0];
  _RAND_1408 = {1{`RANDOM}};
  r_1411 = _RAND_1408[0:0];
  _RAND_1409 = {1{`RANDOM}};
  r_1412 = _RAND_1409[0:0];
  _RAND_1410 = {1{`RANDOM}};
  r_1413 = _RAND_1410[0:0];
  _RAND_1411 = {1{`RANDOM}};
  r_1414 = _RAND_1411[0:0];
  _RAND_1412 = {1{`RANDOM}};
  r_1415 = _RAND_1412[0:0];
  _RAND_1413 = {1{`RANDOM}};
  r_1416 = _RAND_1413[0:0];
  _RAND_1414 = {1{`RANDOM}};
  r_1417 = _RAND_1414[0:0];
  _RAND_1415 = {1{`RANDOM}};
  r_1418 = _RAND_1415[0:0];
  _RAND_1416 = {1{`RANDOM}};
  r_1419 = _RAND_1416[0:0];
  _RAND_1417 = {1{`RANDOM}};
  r_1420 = _RAND_1417[0:0];
  _RAND_1418 = {1{`RANDOM}};
  r_1421 = _RAND_1418[0:0];
  _RAND_1419 = {1{`RANDOM}};
  r_1422 = _RAND_1419[0:0];
  _RAND_1420 = {1{`RANDOM}};
  r_1423 = _RAND_1420[0:0];
  _RAND_1421 = {1{`RANDOM}};
  r_1424 = _RAND_1421[0:0];
  _RAND_1422 = {1{`RANDOM}};
  r_1425 = _RAND_1422[0:0];
  _RAND_1423 = {1{`RANDOM}};
  r_1426 = _RAND_1423[0:0];
  _RAND_1424 = {1{`RANDOM}};
  r_1427 = _RAND_1424[0:0];
  _RAND_1425 = {1{`RANDOM}};
  r_1428 = _RAND_1425[0:0];
  _RAND_1426 = {1{`RANDOM}};
  r_1429 = _RAND_1426[0:0];
  _RAND_1427 = {1{`RANDOM}};
  r_1430 = _RAND_1427[0:0];
  _RAND_1428 = {1{`RANDOM}};
  r_1431 = _RAND_1428[0:0];
  _RAND_1429 = {1{`RANDOM}};
  r_1432 = _RAND_1429[0:0];
  _RAND_1430 = {1{`RANDOM}};
  r_1433 = _RAND_1430[0:0];
  _RAND_1431 = {1{`RANDOM}};
  r_1434 = _RAND_1431[0:0];
  _RAND_1432 = {1{`RANDOM}};
  r_1435 = _RAND_1432[0:0];
  _RAND_1433 = {1{`RANDOM}};
  r_1436 = _RAND_1433[0:0];
  _RAND_1434 = {1{`RANDOM}};
  r_1437 = _RAND_1434[0:0];
  _RAND_1435 = {1{`RANDOM}};
  r_1438 = _RAND_1435[0:0];
  _RAND_1436 = {1{`RANDOM}};
  r_1439 = _RAND_1436[0:0];
  _RAND_1437 = {1{`RANDOM}};
  r_1440 = _RAND_1437[0:0];
  _RAND_1438 = {1{`RANDOM}};
  r_1441 = _RAND_1438[0:0];
  _RAND_1439 = {1{`RANDOM}};
  r_1442 = _RAND_1439[0:0];
  _RAND_1440 = {1{`RANDOM}};
  r_1443 = _RAND_1440[0:0];
  _RAND_1441 = {1{`RANDOM}};
  r_1444 = _RAND_1441[0:0];
  _RAND_1442 = {1{`RANDOM}};
  r_1445 = _RAND_1442[0:0];
  _RAND_1443 = {1{`RANDOM}};
  r_1446 = _RAND_1443[0:0];
  _RAND_1444 = {1{`RANDOM}};
  r_1447 = _RAND_1444[0:0];
  _RAND_1445 = {1{`RANDOM}};
  r_1448 = _RAND_1445[0:0];
  _RAND_1446 = {1{`RANDOM}};
  r_1449 = _RAND_1446[0:0];
  _RAND_1447 = {1{`RANDOM}};
  r_1450 = _RAND_1447[0:0];
  _RAND_1448 = {1{`RANDOM}};
  r_1451 = _RAND_1448[0:0];
  _RAND_1449 = {1{`RANDOM}};
  r_1452 = _RAND_1449[0:0];
  _RAND_1450 = {1{`RANDOM}};
  r_1453 = _RAND_1450[0:0];
  _RAND_1451 = {1{`RANDOM}};
  r_1454 = _RAND_1451[0:0];
  _RAND_1452 = {1{`RANDOM}};
  r_1455 = _RAND_1452[0:0];
  _RAND_1453 = {1{`RANDOM}};
  r_1456 = _RAND_1453[0:0];
  _RAND_1454 = {1{`RANDOM}};
  r_1457 = _RAND_1454[0:0];
  _RAND_1455 = {1{`RANDOM}};
  r_1458 = _RAND_1455[0:0];
  _RAND_1456 = {1{`RANDOM}};
  r_1459 = _RAND_1456[0:0];
  _RAND_1457 = {1{`RANDOM}};
  r_1460 = _RAND_1457[0:0];
  _RAND_1458 = {1{`RANDOM}};
  r_1461 = _RAND_1458[0:0];
  _RAND_1459 = {1{`RANDOM}};
  r_1462 = _RAND_1459[0:0];
  _RAND_1460 = {1{`RANDOM}};
  r_1463 = _RAND_1460[0:0];
  _RAND_1461 = {1{`RANDOM}};
  r_1464 = _RAND_1461[0:0];
  _RAND_1462 = {1{`RANDOM}};
  r_1465 = _RAND_1462[0:0];
  _RAND_1463 = {1{`RANDOM}};
  r_1466 = _RAND_1463[0:0];
  _RAND_1464 = {1{`RANDOM}};
  r_1467 = _RAND_1464[0:0];
  _RAND_1465 = {1{`RANDOM}};
  r_1469 = _RAND_1465[0:0];
  _RAND_1466 = {1{`RANDOM}};
  r_1470 = _RAND_1466[0:0];
  _RAND_1467 = {1{`RANDOM}};
  r_1471 = _RAND_1467[0:0];
  _RAND_1468 = {1{`RANDOM}};
  r_1472 = _RAND_1468[0:0];
  _RAND_1469 = {1{`RANDOM}};
  r_1473 = _RAND_1469[0:0];
  _RAND_1470 = {1{`RANDOM}};
  r_1474 = _RAND_1470[0:0];
  _RAND_1471 = {1{`RANDOM}};
  r_1475 = _RAND_1471[0:0];
  _RAND_1472 = {1{`RANDOM}};
  r_1476 = _RAND_1472[0:0];
  _RAND_1473 = {1{`RANDOM}};
  r_1477 = _RAND_1473[0:0];
  _RAND_1474 = {1{`RANDOM}};
  r_1478 = _RAND_1474[0:0];
  _RAND_1475 = {1{`RANDOM}};
  r_1479 = _RAND_1475[0:0];
  _RAND_1476 = {1{`RANDOM}};
  r_1480 = _RAND_1476[0:0];
  _RAND_1477 = {1{`RANDOM}};
  r_1481 = _RAND_1477[0:0];
  _RAND_1478 = {1{`RANDOM}};
  r_1482 = _RAND_1478[0:0];
  _RAND_1479 = {1{`RANDOM}};
  r_1483 = _RAND_1479[0:0];
  _RAND_1480 = {1{`RANDOM}};
  r_1484 = _RAND_1480[0:0];
  _RAND_1481 = {1{`RANDOM}};
  r_1485 = _RAND_1481[0:0];
  _RAND_1482 = {1{`RANDOM}};
  r_1486 = _RAND_1482[0:0];
  _RAND_1483 = {1{`RANDOM}};
  r_1487 = _RAND_1483[0:0];
  _RAND_1484 = {1{`RANDOM}};
  r_1488 = _RAND_1484[0:0];
  _RAND_1485 = {1{`RANDOM}};
  r_1489 = _RAND_1485[0:0];
  _RAND_1486 = {1{`RANDOM}};
  r_1490 = _RAND_1486[0:0];
  _RAND_1487 = {1{`RANDOM}};
  r_1491 = _RAND_1487[0:0];
  _RAND_1488 = {1{`RANDOM}};
  r_1492 = _RAND_1488[0:0];
  _RAND_1489 = {1{`RANDOM}};
  r_1493 = _RAND_1489[0:0];
  _RAND_1490 = {1{`RANDOM}};
  r_1494 = _RAND_1490[0:0];
  _RAND_1491 = {1{`RANDOM}};
  r_1495 = _RAND_1491[0:0];
  _RAND_1492 = {1{`RANDOM}};
  r_1496 = _RAND_1492[0:0];
  _RAND_1493 = {1{`RANDOM}};
  r_1497 = _RAND_1493[0:0];
  _RAND_1494 = {1{`RANDOM}};
  r_1498 = _RAND_1494[0:0];
  _RAND_1495 = {1{`RANDOM}};
  r_1499 = _RAND_1495[0:0];
  _RAND_1496 = {1{`RANDOM}};
  r_1500 = _RAND_1496[0:0];
  _RAND_1497 = {1{`RANDOM}};
  r_1501 = _RAND_1497[0:0];
  _RAND_1498 = {1{`RANDOM}};
  r_1502 = _RAND_1498[0:0];
  _RAND_1499 = {1{`RANDOM}};
  r_1503 = _RAND_1499[0:0];
  _RAND_1500 = {1{`RANDOM}};
  r_1504 = _RAND_1500[0:0];
  _RAND_1501 = {1{`RANDOM}};
  r_1505 = _RAND_1501[0:0];
  _RAND_1502 = {1{`RANDOM}};
  r_1506 = _RAND_1502[0:0];
  _RAND_1503 = {1{`RANDOM}};
  r_1507 = _RAND_1503[0:0];
  _RAND_1504 = {1{`RANDOM}};
  r_1508 = _RAND_1504[0:0];
  _RAND_1505 = {1{`RANDOM}};
  r_1509 = _RAND_1505[0:0];
  _RAND_1506 = {1{`RANDOM}};
  r_1510 = _RAND_1506[0:0];
  _RAND_1507 = {1{`RANDOM}};
  r_1511 = _RAND_1507[0:0];
  _RAND_1508 = {1{`RANDOM}};
  r_1512 = _RAND_1508[0:0];
  _RAND_1509 = {1{`RANDOM}};
  r_1513 = _RAND_1509[0:0];
  _RAND_1510 = {1{`RANDOM}};
  r_1514 = _RAND_1510[0:0];
  _RAND_1511 = {1{`RANDOM}};
  r_1515 = _RAND_1511[0:0];
  _RAND_1512 = {1{`RANDOM}};
  r_1516 = _RAND_1512[0:0];
  _RAND_1513 = {1{`RANDOM}};
  r_1517 = _RAND_1513[0:0];
  _RAND_1514 = {1{`RANDOM}};
  r_1518 = _RAND_1514[0:0];
  _RAND_1515 = {1{`RANDOM}};
  r_1519 = _RAND_1515[0:0];
  _RAND_1516 = {1{`RANDOM}};
  r_1520 = _RAND_1516[0:0];
  _RAND_1517 = {1{`RANDOM}};
  r_1521 = _RAND_1517[0:0];
  _RAND_1518 = {1{`RANDOM}};
  r_1522 = _RAND_1518[0:0];
  _RAND_1519 = {1{`RANDOM}};
  r_1523 = _RAND_1519[0:0];
  _RAND_1520 = {1{`RANDOM}};
  r_1524 = _RAND_1520[0:0];
  _RAND_1521 = {1{`RANDOM}};
  r_1526 = _RAND_1521[0:0];
  _RAND_1522 = {1{`RANDOM}};
  r_1527 = _RAND_1522[0:0];
  _RAND_1523 = {1{`RANDOM}};
  r_1528 = _RAND_1523[0:0];
  _RAND_1524 = {1{`RANDOM}};
  r_1529 = _RAND_1524[0:0];
  _RAND_1525 = {1{`RANDOM}};
  r_1530 = _RAND_1525[0:0];
  _RAND_1526 = {1{`RANDOM}};
  r_1531 = _RAND_1526[0:0];
  _RAND_1527 = {1{`RANDOM}};
  r_1532 = _RAND_1527[0:0];
  _RAND_1528 = {1{`RANDOM}};
  r_1533 = _RAND_1528[0:0];
  _RAND_1529 = {1{`RANDOM}};
  r_1534 = _RAND_1529[0:0];
  _RAND_1530 = {1{`RANDOM}};
  r_1535 = _RAND_1530[0:0];
  _RAND_1531 = {1{`RANDOM}};
  r_1536 = _RAND_1531[0:0];
  _RAND_1532 = {1{`RANDOM}};
  r_1537 = _RAND_1532[0:0];
  _RAND_1533 = {1{`RANDOM}};
  r_1538 = _RAND_1533[0:0];
  _RAND_1534 = {1{`RANDOM}};
  r_1539 = _RAND_1534[0:0];
  _RAND_1535 = {1{`RANDOM}};
  r_1540 = _RAND_1535[0:0];
  _RAND_1536 = {1{`RANDOM}};
  r_1541 = _RAND_1536[0:0];
  _RAND_1537 = {1{`RANDOM}};
  r_1542 = _RAND_1537[0:0];
  _RAND_1538 = {1{`RANDOM}};
  r_1543 = _RAND_1538[0:0];
  _RAND_1539 = {1{`RANDOM}};
  r_1544 = _RAND_1539[0:0];
  _RAND_1540 = {1{`RANDOM}};
  r_1545 = _RAND_1540[0:0];
  _RAND_1541 = {1{`RANDOM}};
  r_1546 = _RAND_1541[0:0];
  _RAND_1542 = {1{`RANDOM}};
  r_1547 = _RAND_1542[0:0];
  _RAND_1543 = {1{`RANDOM}};
  r_1548 = _RAND_1543[0:0];
  _RAND_1544 = {1{`RANDOM}};
  r_1549 = _RAND_1544[0:0];
  _RAND_1545 = {1{`RANDOM}};
  r_1550 = _RAND_1545[0:0];
  _RAND_1546 = {1{`RANDOM}};
  r_1551 = _RAND_1546[0:0];
  _RAND_1547 = {1{`RANDOM}};
  r_1552 = _RAND_1547[0:0];
  _RAND_1548 = {1{`RANDOM}};
  r_1553 = _RAND_1548[0:0];
  _RAND_1549 = {1{`RANDOM}};
  r_1554 = _RAND_1549[0:0];
  _RAND_1550 = {1{`RANDOM}};
  r_1555 = _RAND_1550[0:0];
  _RAND_1551 = {1{`RANDOM}};
  r_1556 = _RAND_1551[0:0];
  _RAND_1552 = {1{`RANDOM}};
  r_1557 = _RAND_1552[0:0];
  _RAND_1553 = {1{`RANDOM}};
  r_1558 = _RAND_1553[0:0];
  _RAND_1554 = {1{`RANDOM}};
  r_1559 = _RAND_1554[0:0];
  _RAND_1555 = {1{`RANDOM}};
  r_1560 = _RAND_1555[0:0];
  _RAND_1556 = {1{`RANDOM}};
  r_1561 = _RAND_1556[0:0];
  _RAND_1557 = {1{`RANDOM}};
  r_1562 = _RAND_1557[0:0];
  _RAND_1558 = {1{`RANDOM}};
  r_1563 = _RAND_1558[0:0];
  _RAND_1559 = {1{`RANDOM}};
  r_1564 = _RAND_1559[0:0];
  _RAND_1560 = {1{`RANDOM}};
  r_1565 = _RAND_1560[0:0];
  _RAND_1561 = {1{`RANDOM}};
  r_1566 = _RAND_1561[0:0];
  _RAND_1562 = {1{`RANDOM}};
  r_1567 = _RAND_1562[0:0];
  _RAND_1563 = {1{`RANDOM}};
  r_1568 = _RAND_1563[0:0];
  _RAND_1564 = {1{`RANDOM}};
  r_1569 = _RAND_1564[0:0];
  _RAND_1565 = {1{`RANDOM}};
  r_1570 = _RAND_1565[0:0];
  _RAND_1566 = {1{`RANDOM}};
  r_1571 = _RAND_1566[0:0];
  _RAND_1567 = {1{`RANDOM}};
  r_1572 = _RAND_1567[0:0];
  _RAND_1568 = {1{`RANDOM}};
  r_1573 = _RAND_1568[0:0];
  _RAND_1569 = {1{`RANDOM}};
  r_1574 = _RAND_1569[0:0];
  _RAND_1570 = {1{`RANDOM}};
  r_1575 = _RAND_1570[0:0];
  _RAND_1571 = {1{`RANDOM}};
  r_1576 = _RAND_1571[0:0];
  _RAND_1572 = {1{`RANDOM}};
  r_1577 = _RAND_1572[0:0];
  _RAND_1573 = {1{`RANDOM}};
  r_1578 = _RAND_1573[0:0];
  _RAND_1574 = {1{`RANDOM}};
  r_1579 = _RAND_1574[0:0];
  _RAND_1575 = {1{`RANDOM}};
  r_1581 = _RAND_1575[0:0];
  _RAND_1576 = {1{`RANDOM}};
  r_1582 = _RAND_1576[0:0];
  _RAND_1577 = {1{`RANDOM}};
  r_1583 = _RAND_1577[0:0];
  _RAND_1578 = {1{`RANDOM}};
  r_1584 = _RAND_1578[0:0];
  _RAND_1579 = {1{`RANDOM}};
  r_1585 = _RAND_1579[0:0];
  _RAND_1580 = {1{`RANDOM}};
  r_1586 = _RAND_1580[0:0];
  _RAND_1581 = {1{`RANDOM}};
  r_1587 = _RAND_1581[0:0];
  _RAND_1582 = {1{`RANDOM}};
  r_1588 = _RAND_1582[0:0];
  _RAND_1583 = {1{`RANDOM}};
  r_1589 = _RAND_1583[0:0];
  _RAND_1584 = {1{`RANDOM}};
  r_1590 = _RAND_1584[0:0];
  _RAND_1585 = {1{`RANDOM}};
  r_1591 = _RAND_1585[0:0];
  _RAND_1586 = {1{`RANDOM}};
  r_1592 = _RAND_1586[0:0];
  _RAND_1587 = {1{`RANDOM}};
  r_1593 = _RAND_1587[0:0];
  _RAND_1588 = {1{`RANDOM}};
  r_1594 = _RAND_1588[0:0];
  _RAND_1589 = {1{`RANDOM}};
  r_1595 = _RAND_1589[0:0];
  _RAND_1590 = {1{`RANDOM}};
  r_1596 = _RAND_1590[0:0];
  _RAND_1591 = {1{`RANDOM}};
  r_1597 = _RAND_1591[0:0];
  _RAND_1592 = {1{`RANDOM}};
  r_1598 = _RAND_1592[0:0];
  _RAND_1593 = {1{`RANDOM}};
  r_1599 = _RAND_1593[0:0];
  _RAND_1594 = {1{`RANDOM}};
  r_1600 = _RAND_1594[0:0];
  _RAND_1595 = {1{`RANDOM}};
  r_1601 = _RAND_1595[0:0];
  _RAND_1596 = {1{`RANDOM}};
  r_1602 = _RAND_1596[0:0];
  _RAND_1597 = {1{`RANDOM}};
  r_1603 = _RAND_1597[0:0];
  _RAND_1598 = {1{`RANDOM}};
  r_1604 = _RAND_1598[0:0];
  _RAND_1599 = {1{`RANDOM}};
  r_1605 = _RAND_1599[0:0];
  _RAND_1600 = {1{`RANDOM}};
  r_1606 = _RAND_1600[0:0];
  _RAND_1601 = {1{`RANDOM}};
  r_1607 = _RAND_1601[0:0];
  _RAND_1602 = {1{`RANDOM}};
  r_1608 = _RAND_1602[0:0];
  _RAND_1603 = {1{`RANDOM}};
  r_1609 = _RAND_1603[0:0];
  _RAND_1604 = {1{`RANDOM}};
  r_1610 = _RAND_1604[0:0];
  _RAND_1605 = {1{`RANDOM}};
  r_1611 = _RAND_1605[0:0];
  _RAND_1606 = {1{`RANDOM}};
  r_1612 = _RAND_1606[0:0];
  _RAND_1607 = {1{`RANDOM}};
  r_1613 = _RAND_1607[0:0];
  _RAND_1608 = {1{`RANDOM}};
  r_1614 = _RAND_1608[0:0];
  _RAND_1609 = {1{`RANDOM}};
  r_1615 = _RAND_1609[0:0];
  _RAND_1610 = {1{`RANDOM}};
  r_1616 = _RAND_1610[0:0];
  _RAND_1611 = {1{`RANDOM}};
  r_1617 = _RAND_1611[0:0];
  _RAND_1612 = {1{`RANDOM}};
  r_1618 = _RAND_1612[0:0];
  _RAND_1613 = {1{`RANDOM}};
  r_1619 = _RAND_1613[0:0];
  _RAND_1614 = {1{`RANDOM}};
  r_1620 = _RAND_1614[0:0];
  _RAND_1615 = {1{`RANDOM}};
  r_1621 = _RAND_1615[0:0];
  _RAND_1616 = {1{`RANDOM}};
  r_1622 = _RAND_1616[0:0];
  _RAND_1617 = {1{`RANDOM}};
  r_1623 = _RAND_1617[0:0];
  _RAND_1618 = {1{`RANDOM}};
  r_1624 = _RAND_1618[0:0];
  _RAND_1619 = {1{`RANDOM}};
  r_1625 = _RAND_1619[0:0];
  _RAND_1620 = {1{`RANDOM}};
  r_1626 = _RAND_1620[0:0];
  _RAND_1621 = {1{`RANDOM}};
  r_1627 = _RAND_1621[0:0];
  _RAND_1622 = {1{`RANDOM}};
  r_1628 = _RAND_1622[0:0];
  _RAND_1623 = {1{`RANDOM}};
  r_1629 = _RAND_1623[0:0];
  _RAND_1624 = {1{`RANDOM}};
  r_1630 = _RAND_1624[0:0];
  _RAND_1625 = {1{`RANDOM}};
  r_1631 = _RAND_1625[0:0];
  _RAND_1626 = {1{`RANDOM}};
  r_1632 = _RAND_1626[0:0];
  _RAND_1627 = {1{`RANDOM}};
  r_1634 = _RAND_1627[0:0];
  _RAND_1628 = {1{`RANDOM}};
  r_1635 = _RAND_1628[0:0];
  _RAND_1629 = {1{`RANDOM}};
  r_1636 = _RAND_1629[0:0];
  _RAND_1630 = {1{`RANDOM}};
  r_1637 = _RAND_1630[0:0];
  _RAND_1631 = {1{`RANDOM}};
  r_1638 = _RAND_1631[0:0];
  _RAND_1632 = {1{`RANDOM}};
  r_1639 = _RAND_1632[0:0];
  _RAND_1633 = {1{`RANDOM}};
  r_1640 = _RAND_1633[0:0];
  _RAND_1634 = {1{`RANDOM}};
  r_1641 = _RAND_1634[0:0];
  _RAND_1635 = {1{`RANDOM}};
  r_1642 = _RAND_1635[0:0];
  _RAND_1636 = {1{`RANDOM}};
  r_1643 = _RAND_1636[0:0];
  _RAND_1637 = {1{`RANDOM}};
  r_1644 = _RAND_1637[0:0];
  _RAND_1638 = {1{`RANDOM}};
  r_1645 = _RAND_1638[0:0];
  _RAND_1639 = {1{`RANDOM}};
  r_1646 = _RAND_1639[0:0];
  _RAND_1640 = {1{`RANDOM}};
  r_1647 = _RAND_1640[0:0];
  _RAND_1641 = {1{`RANDOM}};
  r_1648 = _RAND_1641[0:0];
  _RAND_1642 = {1{`RANDOM}};
  r_1649 = _RAND_1642[0:0];
  _RAND_1643 = {1{`RANDOM}};
  r_1650 = _RAND_1643[0:0];
  _RAND_1644 = {1{`RANDOM}};
  r_1651 = _RAND_1644[0:0];
  _RAND_1645 = {1{`RANDOM}};
  r_1652 = _RAND_1645[0:0];
  _RAND_1646 = {1{`RANDOM}};
  r_1653 = _RAND_1646[0:0];
  _RAND_1647 = {1{`RANDOM}};
  r_1654 = _RAND_1647[0:0];
  _RAND_1648 = {1{`RANDOM}};
  r_1655 = _RAND_1648[0:0];
  _RAND_1649 = {1{`RANDOM}};
  r_1656 = _RAND_1649[0:0];
  _RAND_1650 = {1{`RANDOM}};
  r_1657 = _RAND_1650[0:0];
  _RAND_1651 = {1{`RANDOM}};
  r_1658 = _RAND_1651[0:0];
  _RAND_1652 = {1{`RANDOM}};
  r_1659 = _RAND_1652[0:0];
  _RAND_1653 = {1{`RANDOM}};
  r_1660 = _RAND_1653[0:0];
  _RAND_1654 = {1{`RANDOM}};
  r_1661 = _RAND_1654[0:0];
  _RAND_1655 = {1{`RANDOM}};
  r_1662 = _RAND_1655[0:0];
  _RAND_1656 = {1{`RANDOM}};
  r_1663 = _RAND_1656[0:0];
  _RAND_1657 = {1{`RANDOM}};
  r_1664 = _RAND_1657[0:0];
  _RAND_1658 = {1{`RANDOM}};
  r_1665 = _RAND_1658[0:0];
  _RAND_1659 = {1{`RANDOM}};
  r_1666 = _RAND_1659[0:0];
  _RAND_1660 = {1{`RANDOM}};
  r_1667 = _RAND_1660[0:0];
  _RAND_1661 = {1{`RANDOM}};
  r_1668 = _RAND_1661[0:0];
  _RAND_1662 = {1{`RANDOM}};
  r_1669 = _RAND_1662[0:0];
  _RAND_1663 = {1{`RANDOM}};
  r_1670 = _RAND_1663[0:0];
  _RAND_1664 = {1{`RANDOM}};
  r_1671 = _RAND_1664[0:0];
  _RAND_1665 = {1{`RANDOM}};
  r_1672 = _RAND_1665[0:0];
  _RAND_1666 = {1{`RANDOM}};
  r_1673 = _RAND_1666[0:0];
  _RAND_1667 = {1{`RANDOM}};
  r_1674 = _RAND_1667[0:0];
  _RAND_1668 = {1{`RANDOM}};
  r_1675 = _RAND_1668[0:0];
  _RAND_1669 = {1{`RANDOM}};
  r_1676 = _RAND_1669[0:0];
  _RAND_1670 = {1{`RANDOM}};
  r_1677 = _RAND_1670[0:0];
  _RAND_1671 = {1{`RANDOM}};
  r_1678 = _RAND_1671[0:0];
  _RAND_1672 = {1{`RANDOM}};
  r_1679 = _RAND_1672[0:0];
  _RAND_1673 = {1{`RANDOM}};
  r_1680 = _RAND_1673[0:0];
  _RAND_1674 = {1{`RANDOM}};
  r_1681 = _RAND_1674[0:0];
  _RAND_1675 = {1{`RANDOM}};
  r_1682 = _RAND_1675[0:0];
  _RAND_1676 = {1{`RANDOM}};
  r_1683 = _RAND_1676[0:0];
  _RAND_1677 = {1{`RANDOM}};
  r_1685 = _RAND_1677[0:0];
  _RAND_1678 = {1{`RANDOM}};
  r_1686 = _RAND_1678[0:0];
  _RAND_1679 = {1{`RANDOM}};
  r_1687 = _RAND_1679[0:0];
  _RAND_1680 = {1{`RANDOM}};
  r_1688 = _RAND_1680[0:0];
  _RAND_1681 = {1{`RANDOM}};
  r_1689 = _RAND_1681[0:0];
  _RAND_1682 = {1{`RANDOM}};
  r_1690 = _RAND_1682[0:0];
  _RAND_1683 = {1{`RANDOM}};
  r_1691 = _RAND_1683[0:0];
  _RAND_1684 = {1{`RANDOM}};
  r_1692 = _RAND_1684[0:0];
  _RAND_1685 = {1{`RANDOM}};
  r_1693 = _RAND_1685[0:0];
  _RAND_1686 = {1{`RANDOM}};
  r_1694 = _RAND_1686[0:0];
  _RAND_1687 = {1{`RANDOM}};
  r_1695 = _RAND_1687[0:0];
  _RAND_1688 = {1{`RANDOM}};
  r_1696 = _RAND_1688[0:0];
  _RAND_1689 = {1{`RANDOM}};
  r_1697 = _RAND_1689[0:0];
  _RAND_1690 = {1{`RANDOM}};
  r_1698 = _RAND_1690[0:0];
  _RAND_1691 = {1{`RANDOM}};
  r_1699 = _RAND_1691[0:0];
  _RAND_1692 = {1{`RANDOM}};
  r_1700 = _RAND_1692[0:0];
  _RAND_1693 = {1{`RANDOM}};
  r_1701 = _RAND_1693[0:0];
  _RAND_1694 = {1{`RANDOM}};
  r_1702 = _RAND_1694[0:0];
  _RAND_1695 = {1{`RANDOM}};
  r_1703 = _RAND_1695[0:0];
  _RAND_1696 = {1{`RANDOM}};
  r_1704 = _RAND_1696[0:0];
  _RAND_1697 = {1{`RANDOM}};
  r_1705 = _RAND_1697[0:0];
  _RAND_1698 = {1{`RANDOM}};
  r_1706 = _RAND_1698[0:0];
  _RAND_1699 = {1{`RANDOM}};
  r_1707 = _RAND_1699[0:0];
  _RAND_1700 = {1{`RANDOM}};
  r_1708 = _RAND_1700[0:0];
  _RAND_1701 = {1{`RANDOM}};
  r_1709 = _RAND_1701[0:0];
  _RAND_1702 = {1{`RANDOM}};
  r_1710 = _RAND_1702[0:0];
  _RAND_1703 = {1{`RANDOM}};
  r_1711 = _RAND_1703[0:0];
  _RAND_1704 = {1{`RANDOM}};
  r_1712 = _RAND_1704[0:0];
  _RAND_1705 = {1{`RANDOM}};
  r_1713 = _RAND_1705[0:0];
  _RAND_1706 = {1{`RANDOM}};
  r_1714 = _RAND_1706[0:0];
  _RAND_1707 = {1{`RANDOM}};
  r_1715 = _RAND_1707[0:0];
  _RAND_1708 = {1{`RANDOM}};
  r_1716 = _RAND_1708[0:0];
  _RAND_1709 = {1{`RANDOM}};
  r_1717 = _RAND_1709[0:0];
  _RAND_1710 = {1{`RANDOM}};
  r_1718 = _RAND_1710[0:0];
  _RAND_1711 = {1{`RANDOM}};
  r_1719 = _RAND_1711[0:0];
  _RAND_1712 = {1{`RANDOM}};
  r_1720 = _RAND_1712[0:0];
  _RAND_1713 = {1{`RANDOM}};
  r_1721 = _RAND_1713[0:0];
  _RAND_1714 = {1{`RANDOM}};
  r_1722 = _RAND_1714[0:0];
  _RAND_1715 = {1{`RANDOM}};
  r_1723 = _RAND_1715[0:0];
  _RAND_1716 = {1{`RANDOM}};
  r_1724 = _RAND_1716[0:0];
  _RAND_1717 = {1{`RANDOM}};
  r_1725 = _RAND_1717[0:0];
  _RAND_1718 = {1{`RANDOM}};
  r_1726 = _RAND_1718[0:0];
  _RAND_1719 = {1{`RANDOM}};
  r_1727 = _RAND_1719[0:0];
  _RAND_1720 = {1{`RANDOM}};
  r_1728 = _RAND_1720[0:0];
  _RAND_1721 = {1{`RANDOM}};
  r_1729 = _RAND_1721[0:0];
  _RAND_1722 = {1{`RANDOM}};
  r_1730 = _RAND_1722[0:0];
  _RAND_1723 = {1{`RANDOM}};
  r_1731 = _RAND_1723[0:0];
  _RAND_1724 = {1{`RANDOM}};
  r_1732 = _RAND_1724[0:0];
  _RAND_1725 = {1{`RANDOM}};
  r_1734 = _RAND_1725[0:0];
  _RAND_1726 = {1{`RANDOM}};
  r_1735 = _RAND_1726[0:0];
  _RAND_1727 = {1{`RANDOM}};
  r_1736 = _RAND_1727[0:0];
  _RAND_1728 = {1{`RANDOM}};
  r_1737 = _RAND_1728[0:0];
  _RAND_1729 = {1{`RANDOM}};
  r_1738 = _RAND_1729[0:0];
  _RAND_1730 = {1{`RANDOM}};
  r_1739 = _RAND_1730[0:0];
  _RAND_1731 = {1{`RANDOM}};
  r_1740 = _RAND_1731[0:0];
  _RAND_1732 = {1{`RANDOM}};
  r_1741 = _RAND_1732[0:0];
  _RAND_1733 = {1{`RANDOM}};
  r_1742 = _RAND_1733[0:0];
  _RAND_1734 = {1{`RANDOM}};
  r_1743 = _RAND_1734[0:0];
  _RAND_1735 = {1{`RANDOM}};
  r_1744 = _RAND_1735[0:0];
  _RAND_1736 = {1{`RANDOM}};
  r_1745 = _RAND_1736[0:0];
  _RAND_1737 = {1{`RANDOM}};
  r_1746 = _RAND_1737[0:0];
  _RAND_1738 = {1{`RANDOM}};
  r_1747 = _RAND_1738[0:0];
  _RAND_1739 = {1{`RANDOM}};
  r_1748 = _RAND_1739[0:0];
  _RAND_1740 = {1{`RANDOM}};
  r_1749 = _RAND_1740[0:0];
  _RAND_1741 = {1{`RANDOM}};
  r_1750 = _RAND_1741[0:0];
  _RAND_1742 = {1{`RANDOM}};
  r_1751 = _RAND_1742[0:0];
  _RAND_1743 = {1{`RANDOM}};
  r_1752 = _RAND_1743[0:0];
  _RAND_1744 = {1{`RANDOM}};
  r_1753 = _RAND_1744[0:0];
  _RAND_1745 = {1{`RANDOM}};
  r_1754 = _RAND_1745[0:0];
  _RAND_1746 = {1{`RANDOM}};
  r_1755 = _RAND_1746[0:0];
  _RAND_1747 = {1{`RANDOM}};
  r_1756 = _RAND_1747[0:0];
  _RAND_1748 = {1{`RANDOM}};
  r_1757 = _RAND_1748[0:0];
  _RAND_1749 = {1{`RANDOM}};
  r_1758 = _RAND_1749[0:0];
  _RAND_1750 = {1{`RANDOM}};
  r_1759 = _RAND_1750[0:0];
  _RAND_1751 = {1{`RANDOM}};
  r_1760 = _RAND_1751[0:0];
  _RAND_1752 = {1{`RANDOM}};
  r_1761 = _RAND_1752[0:0];
  _RAND_1753 = {1{`RANDOM}};
  r_1762 = _RAND_1753[0:0];
  _RAND_1754 = {1{`RANDOM}};
  r_1763 = _RAND_1754[0:0];
  _RAND_1755 = {1{`RANDOM}};
  r_1764 = _RAND_1755[0:0];
  _RAND_1756 = {1{`RANDOM}};
  r_1765 = _RAND_1756[0:0];
  _RAND_1757 = {1{`RANDOM}};
  r_1766 = _RAND_1757[0:0];
  _RAND_1758 = {1{`RANDOM}};
  r_1767 = _RAND_1758[0:0];
  _RAND_1759 = {1{`RANDOM}};
  r_1768 = _RAND_1759[0:0];
  _RAND_1760 = {1{`RANDOM}};
  r_1769 = _RAND_1760[0:0];
  _RAND_1761 = {1{`RANDOM}};
  r_1770 = _RAND_1761[0:0];
  _RAND_1762 = {1{`RANDOM}};
  r_1771 = _RAND_1762[0:0];
  _RAND_1763 = {1{`RANDOM}};
  r_1772 = _RAND_1763[0:0];
  _RAND_1764 = {1{`RANDOM}};
  r_1773 = _RAND_1764[0:0];
  _RAND_1765 = {1{`RANDOM}};
  r_1774 = _RAND_1765[0:0];
  _RAND_1766 = {1{`RANDOM}};
  r_1775 = _RAND_1766[0:0];
  _RAND_1767 = {1{`RANDOM}};
  r_1776 = _RAND_1767[0:0];
  _RAND_1768 = {1{`RANDOM}};
  r_1777 = _RAND_1768[0:0];
  _RAND_1769 = {1{`RANDOM}};
  r_1778 = _RAND_1769[0:0];
  _RAND_1770 = {1{`RANDOM}};
  r_1779 = _RAND_1770[0:0];
  _RAND_1771 = {1{`RANDOM}};
  r_1781 = _RAND_1771[0:0];
  _RAND_1772 = {1{`RANDOM}};
  r_1782 = _RAND_1772[0:0];
  _RAND_1773 = {1{`RANDOM}};
  r_1783 = _RAND_1773[0:0];
  _RAND_1774 = {1{`RANDOM}};
  r_1784 = _RAND_1774[0:0];
  _RAND_1775 = {1{`RANDOM}};
  r_1785 = _RAND_1775[0:0];
  _RAND_1776 = {1{`RANDOM}};
  r_1786 = _RAND_1776[0:0];
  _RAND_1777 = {1{`RANDOM}};
  r_1787 = _RAND_1777[0:0];
  _RAND_1778 = {1{`RANDOM}};
  r_1788 = _RAND_1778[0:0];
  _RAND_1779 = {1{`RANDOM}};
  r_1789 = _RAND_1779[0:0];
  _RAND_1780 = {1{`RANDOM}};
  r_1790 = _RAND_1780[0:0];
  _RAND_1781 = {1{`RANDOM}};
  r_1791 = _RAND_1781[0:0];
  _RAND_1782 = {1{`RANDOM}};
  r_1792 = _RAND_1782[0:0];
  _RAND_1783 = {1{`RANDOM}};
  r_1793 = _RAND_1783[0:0];
  _RAND_1784 = {1{`RANDOM}};
  r_1794 = _RAND_1784[0:0];
  _RAND_1785 = {1{`RANDOM}};
  r_1795 = _RAND_1785[0:0];
  _RAND_1786 = {1{`RANDOM}};
  r_1796 = _RAND_1786[0:0];
  _RAND_1787 = {1{`RANDOM}};
  r_1797 = _RAND_1787[0:0];
  _RAND_1788 = {1{`RANDOM}};
  r_1798 = _RAND_1788[0:0];
  _RAND_1789 = {1{`RANDOM}};
  r_1799 = _RAND_1789[0:0];
  _RAND_1790 = {1{`RANDOM}};
  r_1800 = _RAND_1790[0:0];
  _RAND_1791 = {1{`RANDOM}};
  r_1801 = _RAND_1791[0:0];
  _RAND_1792 = {1{`RANDOM}};
  r_1802 = _RAND_1792[0:0];
  _RAND_1793 = {1{`RANDOM}};
  r_1803 = _RAND_1793[0:0];
  _RAND_1794 = {1{`RANDOM}};
  r_1804 = _RAND_1794[0:0];
  _RAND_1795 = {1{`RANDOM}};
  r_1805 = _RAND_1795[0:0];
  _RAND_1796 = {1{`RANDOM}};
  r_1806 = _RAND_1796[0:0];
  _RAND_1797 = {1{`RANDOM}};
  r_1807 = _RAND_1797[0:0];
  _RAND_1798 = {1{`RANDOM}};
  r_1808 = _RAND_1798[0:0];
  _RAND_1799 = {1{`RANDOM}};
  r_1809 = _RAND_1799[0:0];
  _RAND_1800 = {1{`RANDOM}};
  r_1810 = _RAND_1800[0:0];
  _RAND_1801 = {1{`RANDOM}};
  r_1811 = _RAND_1801[0:0];
  _RAND_1802 = {1{`RANDOM}};
  r_1812 = _RAND_1802[0:0];
  _RAND_1803 = {1{`RANDOM}};
  r_1813 = _RAND_1803[0:0];
  _RAND_1804 = {1{`RANDOM}};
  r_1814 = _RAND_1804[0:0];
  _RAND_1805 = {1{`RANDOM}};
  r_1815 = _RAND_1805[0:0];
  _RAND_1806 = {1{`RANDOM}};
  r_1816 = _RAND_1806[0:0];
  _RAND_1807 = {1{`RANDOM}};
  r_1817 = _RAND_1807[0:0];
  _RAND_1808 = {1{`RANDOM}};
  r_1818 = _RAND_1808[0:0];
  _RAND_1809 = {1{`RANDOM}};
  r_1819 = _RAND_1809[0:0];
  _RAND_1810 = {1{`RANDOM}};
  r_1820 = _RAND_1810[0:0];
  _RAND_1811 = {1{`RANDOM}};
  r_1821 = _RAND_1811[0:0];
  _RAND_1812 = {1{`RANDOM}};
  r_1822 = _RAND_1812[0:0];
  _RAND_1813 = {1{`RANDOM}};
  r_1823 = _RAND_1813[0:0];
  _RAND_1814 = {1{`RANDOM}};
  r_1824 = _RAND_1814[0:0];
  _RAND_1815 = {1{`RANDOM}};
  r_1826 = _RAND_1815[0:0];
  _RAND_1816 = {1{`RANDOM}};
  r_1827 = _RAND_1816[0:0];
  _RAND_1817 = {1{`RANDOM}};
  r_1828 = _RAND_1817[0:0];
  _RAND_1818 = {1{`RANDOM}};
  r_1829 = _RAND_1818[0:0];
  _RAND_1819 = {1{`RANDOM}};
  r_1830 = _RAND_1819[0:0];
  _RAND_1820 = {1{`RANDOM}};
  r_1831 = _RAND_1820[0:0];
  _RAND_1821 = {1{`RANDOM}};
  r_1832 = _RAND_1821[0:0];
  _RAND_1822 = {1{`RANDOM}};
  r_1833 = _RAND_1822[0:0];
  _RAND_1823 = {1{`RANDOM}};
  r_1834 = _RAND_1823[0:0];
  _RAND_1824 = {1{`RANDOM}};
  r_1835 = _RAND_1824[0:0];
  _RAND_1825 = {1{`RANDOM}};
  r_1836 = _RAND_1825[0:0];
  _RAND_1826 = {1{`RANDOM}};
  r_1837 = _RAND_1826[0:0];
  _RAND_1827 = {1{`RANDOM}};
  r_1838 = _RAND_1827[0:0];
  _RAND_1828 = {1{`RANDOM}};
  r_1839 = _RAND_1828[0:0];
  _RAND_1829 = {1{`RANDOM}};
  r_1840 = _RAND_1829[0:0];
  _RAND_1830 = {1{`RANDOM}};
  r_1841 = _RAND_1830[0:0];
  _RAND_1831 = {1{`RANDOM}};
  r_1842 = _RAND_1831[0:0];
  _RAND_1832 = {1{`RANDOM}};
  r_1843 = _RAND_1832[0:0];
  _RAND_1833 = {1{`RANDOM}};
  r_1844 = _RAND_1833[0:0];
  _RAND_1834 = {1{`RANDOM}};
  r_1845 = _RAND_1834[0:0];
  _RAND_1835 = {1{`RANDOM}};
  r_1846 = _RAND_1835[0:0];
  _RAND_1836 = {1{`RANDOM}};
  r_1847 = _RAND_1836[0:0];
  _RAND_1837 = {1{`RANDOM}};
  r_1848 = _RAND_1837[0:0];
  _RAND_1838 = {1{`RANDOM}};
  r_1849 = _RAND_1838[0:0];
  _RAND_1839 = {1{`RANDOM}};
  r_1850 = _RAND_1839[0:0];
  _RAND_1840 = {1{`RANDOM}};
  r_1851 = _RAND_1840[0:0];
  _RAND_1841 = {1{`RANDOM}};
  r_1852 = _RAND_1841[0:0];
  _RAND_1842 = {1{`RANDOM}};
  r_1853 = _RAND_1842[0:0];
  _RAND_1843 = {1{`RANDOM}};
  r_1854 = _RAND_1843[0:0];
  _RAND_1844 = {1{`RANDOM}};
  r_1855 = _RAND_1844[0:0];
  _RAND_1845 = {1{`RANDOM}};
  r_1856 = _RAND_1845[0:0];
  _RAND_1846 = {1{`RANDOM}};
  r_1857 = _RAND_1846[0:0];
  _RAND_1847 = {1{`RANDOM}};
  r_1858 = _RAND_1847[0:0];
  _RAND_1848 = {1{`RANDOM}};
  r_1859 = _RAND_1848[0:0];
  _RAND_1849 = {1{`RANDOM}};
  r_1860 = _RAND_1849[0:0];
  _RAND_1850 = {1{`RANDOM}};
  r_1861 = _RAND_1850[0:0];
  _RAND_1851 = {1{`RANDOM}};
  r_1862 = _RAND_1851[0:0];
  _RAND_1852 = {1{`RANDOM}};
  r_1863 = _RAND_1852[0:0];
  _RAND_1853 = {1{`RANDOM}};
  r_1864 = _RAND_1853[0:0];
  _RAND_1854 = {1{`RANDOM}};
  r_1865 = _RAND_1854[0:0];
  _RAND_1855 = {1{`RANDOM}};
  r_1866 = _RAND_1855[0:0];
  _RAND_1856 = {1{`RANDOM}};
  r_1867 = _RAND_1856[0:0];
  _RAND_1857 = {1{`RANDOM}};
  r_1869 = _RAND_1857[0:0];
  _RAND_1858 = {1{`RANDOM}};
  r_1870 = _RAND_1858[0:0];
  _RAND_1859 = {1{`RANDOM}};
  r_1871 = _RAND_1859[0:0];
  _RAND_1860 = {1{`RANDOM}};
  r_1872 = _RAND_1860[0:0];
  _RAND_1861 = {1{`RANDOM}};
  r_1873 = _RAND_1861[0:0];
  _RAND_1862 = {1{`RANDOM}};
  r_1874 = _RAND_1862[0:0];
  _RAND_1863 = {1{`RANDOM}};
  r_1875 = _RAND_1863[0:0];
  _RAND_1864 = {1{`RANDOM}};
  r_1876 = _RAND_1864[0:0];
  _RAND_1865 = {1{`RANDOM}};
  r_1877 = _RAND_1865[0:0];
  _RAND_1866 = {1{`RANDOM}};
  r_1878 = _RAND_1866[0:0];
  _RAND_1867 = {1{`RANDOM}};
  r_1879 = _RAND_1867[0:0];
  _RAND_1868 = {1{`RANDOM}};
  r_1880 = _RAND_1868[0:0];
  _RAND_1869 = {1{`RANDOM}};
  r_1881 = _RAND_1869[0:0];
  _RAND_1870 = {1{`RANDOM}};
  r_1882 = _RAND_1870[0:0];
  _RAND_1871 = {1{`RANDOM}};
  r_1883 = _RAND_1871[0:0];
  _RAND_1872 = {1{`RANDOM}};
  r_1884 = _RAND_1872[0:0];
  _RAND_1873 = {1{`RANDOM}};
  r_1885 = _RAND_1873[0:0];
  _RAND_1874 = {1{`RANDOM}};
  r_1886 = _RAND_1874[0:0];
  _RAND_1875 = {1{`RANDOM}};
  r_1887 = _RAND_1875[0:0];
  _RAND_1876 = {1{`RANDOM}};
  r_1888 = _RAND_1876[0:0];
  _RAND_1877 = {1{`RANDOM}};
  r_1889 = _RAND_1877[0:0];
  _RAND_1878 = {1{`RANDOM}};
  r_1890 = _RAND_1878[0:0];
  _RAND_1879 = {1{`RANDOM}};
  r_1891 = _RAND_1879[0:0];
  _RAND_1880 = {1{`RANDOM}};
  r_1892 = _RAND_1880[0:0];
  _RAND_1881 = {1{`RANDOM}};
  r_1893 = _RAND_1881[0:0];
  _RAND_1882 = {1{`RANDOM}};
  r_1894 = _RAND_1882[0:0];
  _RAND_1883 = {1{`RANDOM}};
  r_1895 = _RAND_1883[0:0];
  _RAND_1884 = {1{`RANDOM}};
  r_1896 = _RAND_1884[0:0];
  _RAND_1885 = {1{`RANDOM}};
  r_1897 = _RAND_1885[0:0];
  _RAND_1886 = {1{`RANDOM}};
  r_1898 = _RAND_1886[0:0];
  _RAND_1887 = {1{`RANDOM}};
  r_1899 = _RAND_1887[0:0];
  _RAND_1888 = {1{`RANDOM}};
  r_1900 = _RAND_1888[0:0];
  _RAND_1889 = {1{`RANDOM}};
  r_1901 = _RAND_1889[0:0];
  _RAND_1890 = {1{`RANDOM}};
  r_1902 = _RAND_1890[0:0];
  _RAND_1891 = {1{`RANDOM}};
  r_1903 = _RAND_1891[0:0];
  _RAND_1892 = {1{`RANDOM}};
  r_1904 = _RAND_1892[0:0];
  _RAND_1893 = {1{`RANDOM}};
  r_1905 = _RAND_1893[0:0];
  _RAND_1894 = {1{`RANDOM}};
  r_1906 = _RAND_1894[0:0];
  _RAND_1895 = {1{`RANDOM}};
  r_1907 = _RAND_1895[0:0];
  _RAND_1896 = {1{`RANDOM}};
  r_1908 = _RAND_1896[0:0];
  _RAND_1897 = {1{`RANDOM}};
  r_1910 = _RAND_1897[0:0];
  _RAND_1898 = {1{`RANDOM}};
  r_1911 = _RAND_1898[0:0];
  _RAND_1899 = {1{`RANDOM}};
  r_1912 = _RAND_1899[0:0];
  _RAND_1900 = {1{`RANDOM}};
  r_1913 = _RAND_1900[0:0];
  _RAND_1901 = {1{`RANDOM}};
  r_1914 = _RAND_1901[0:0];
  _RAND_1902 = {1{`RANDOM}};
  r_1915 = _RAND_1902[0:0];
  _RAND_1903 = {1{`RANDOM}};
  r_1916 = _RAND_1903[0:0];
  _RAND_1904 = {1{`RANDOM}};
  r_1917 = _RAND_1904[0:0];
  _RAND_1905 = {1{`RANDOM}};
  r_1918 = _RAND_1905[0:0];
  _RAND_1906 = {1{`RANDOM}};
  r_1919 = _RAND_1906[0:0];
  _RAND_1907 = {1{`RANDOM}};
  r_1920 = _RAND_1907[0:0];
  _RAND_1908 = {1{`RANDOM}};
  r_1921 = _RAND_1908[0:0];
  _RAND_1909 = {1{`RANDOM}};
  r_1922 = _RAND_1909[0:0];
  _RAND_1910 = {1{`RANDOM}};
  r_1923 = _RAND_1910[0:0];
  _RAND_1911 = {1{`RANDOM}};
  r_1924 = _RAND_1911[0:0];
  _RAND_1912 = {1{`RANDOM}};
  r_1925 = _RAND_1912[0:0];
  _RAND_1913 = {1{`RANDOM}};
  r_1926 = _RAND_1913[0:0];
  _RAND_1914 = {1{`RANDOM}};
  r_1927 = _RAND_1914[0:0];
  _RAND_1915 = {1{`RANDOM}};
  r_1928 = _RAND_1915[0:0];
  _RAND_1916 = {1{`RANDOM}};
  r_1929 = _RAND_1916[0:0];
  _RAND_1917 = {1{`RANDOM}};
  r_1930 = _RAND_1917[0:0];
  _RAND_1918 = {1{`RANDOM}};
  r_1931 = _RAND_1918[0:0];
  _RAND_1919 = {1{`RANDOM}};
  r_1932 = _RAND_1919[0:0];
  _RAND_1920 = {1{`RANDOM}};
  r_1933 = _RAND_1920[0:0];
  _RAND_1921 = {1{`RANDOM}};
  r_1934 = _RAND_1921[0:0];
  _RAND_1922 = {1{`RANDOM}};
  r_1935 = _RAND_1922[0:0];
  _RAND_1923 = {1{`RANDOM}};
  r_1936 = _RAND_1923[0:0];
  _RAND_1924 = {1{`RANDOM}};
  r_1937 = _RAND_1924[0:0];
  _RAND_1925 = {1{`RANDOM}};
  r_1938 = _RAND_1925[0:0];
  _RAND_1926 = {1{`RANDOM}};
  r_1939 = _RAND_1926[0:0];
  _RAND_1927 = {1{`RANDOM}};
  r_1940 = _RAND_1927[0:0];
  _RAND_1928 = {1{`RANDOM}};
  r_1941 = _RAND_1928[0:0];
  _RAND_1929 = {1{`RANDOM}};
  r_1942 = _RAND_1929[0:0];
  _RAND_1930 = {1{`RANDOM}};
  r_1943 = _RAND_1930[0:0];
  _RAND_1931 = {1{`RANDOM}};
  r_1944 = _RAND_1931[0:0];
  _RAND_1932 = {1{`RANDOM}};
  r_1945 = _RAND_1932[0:0];
  _RAND_1933 = {1{`RANDOM}};
  r_1946 = _RAND_1933[0:0];
  _RAND_1934 = {1{`RANDOM}};
  r_1947 = _RAND_1934[0:0];
  _RAND_1935 = {1{`RANDOM}};
  r_1949 = _RAND_1935[0:0];
  _RAND_1936 = {1{`RANDOM}};
  r_1950 = _RAND_1936[0:0];
  _RAND_1937 = {1{`RANDOM}};
  r_1951 = _RAND_1937[0:0];
  _RAND_1938 = {1{`RANDOM}};
  r_1952 = _RAND_1938[0:0];
  _RAND_1939 = {1{`RANDOM}};
  r_1953 = _RAND_1939[0:0];
  _RAND_1940 = {1{`RANDOM}};
  r_1954 = _RAND_1940[0:0];
  _RAND_1941 = {1{`RANDOM}};
  r_1955 = _RAND_1941[0:0];
  _RAND_1942 = {1{`RANDOM}};
  r_1956 = _RAND_1942[0:0];
  _RAND_1943 = {1{`RANDOM}};
  r_1957 = _RAND_1943[0:0];
  _RAND_1944 = {1{`RANDOM}};
  r_1958 = _RAND_1944[0:0];
  _RAND_1945 = {1{`RANDOM}};
  r_1959 = _RAND_1945[0:0];
  _RAND_1946 = {1{`RANDOM}};
  r_1960 = _RAND_1946[0:0];
  _RAND_1947 = {1{`RANDOM}};
  r_1961 = _RAND_1947[0:0];
  _RAND_1948 = {1{`RANDOM}};
  r_1962 = _RAND_1948[0:0];
  _RAND_1949 = {1{`RANDOM}};
  r_1963 = _RAND_1949[0:0];
  _RAND_1950 = {1{`RANDOM}};
  r_1964 = _RAND_1950[0:0];
  _RAND_1951 = {1{`RANDOM}};
  r_1965 = _RAND_1951[0:0];
  _RAND_1952 = {1{`RANDOM}};
  r_1966 = _RAND_1952[0:0];
  _RAND_1953 = {1{`RANDOM}};
  r_1967 = _RAND_1953[0:0];
  _RAND_1954 = {1{`RANDOM}};
  r_1968 = _RAND_1954[0:0];
  _RAND_1955 = {1{`RANDOM}};
  r_1969 = _RAND_1955[0:0];
  _RAND_1956 = {1{`RANDOM}};
  r_1970 = _RAND_1956[0:0];
  _RAND_1957 = {1{`RANDOM}};
  r_1971 = _RAND_1957[0:0];
  _RAND_1958 = {1{`RANDOM}};
  r_1972 = _RAND_1958[0:0];
  _RAND_1959 = {1{`RANDOM}};
  r_1973 = _RAND_1959[0:0];
  _RAND_1960 = {1{`RANDOM}};
  r_1974 = _RAND_1960[0:0];
  _RAND_1961 = {1{`RANDOM}};
  r_1975 = _RAND_1961[0:0];
  _RAND_1962 = {1{`RANDOM}};
  r_1976 = _RAND_1962[0:0];
  _RAND_1963 = {1{`RANDOM}};
  r_1977 = _RAND_1963[0:0];
  _RAND_1964 = {1{`RANDOM}};
  r_1978 = _RAND_1964[0:0];
  _RAND_1965 = {1{`RANDOM}};
  r_1979 = _RAND_1965[0:0];
  _RAND_1966 = {1{`RANDOM}};
  r_1980 = _RAND_1966[0:0];
  _RAND_1967 = {1{`RANDOM}};
  r_1981 = _RAND_1967[0:0];
  _RAND_1968 = {1{`RANDOM}};
  r_1982 = _RAND_1968[0:0];
  _RAND_1969 = {1{`RANDOM}};
  r_1983 = _RAND_1969[0:0];
  _RAND_1970 = {1{`RANDOM}};
  r_1984 = _RAND_1970[0:0];
  _RAND_1971 = {1{`RANDOM}};
  r_1986 = _RAND_1971[0:0];
  _RAND_1972 = {1{`RANDOM}};
  r_1987 = _RAND_1972[0:0];
  _RAND_1973 = {1{`RANDOM}};
  r_1988 = _RAND_1973[0:0];
  _RAND_1974 = {1{`RANDOM}};
  r_1989 = _RAND_1974[0:0];
  _RAND_1975 = {1{`RANDOM}};
  r_1990 = _RAND_1975[0:0];
  _RAND_1976 = {1{`RANDOM}};
  r_1991 = _RAND_1976[0:0];
  _RAND_1977 = {1{`RANDOM}};
  r_1992 = _RAND_1977[0:0];
  _RAND_1978 = {1{`RANDOM}};
  r_1993 = _RAND_1978[0:0];
  _RAND_1979 = {1{`RANDOM}};
  r_1994 = _RAND_1979[0:0];
  _RAND_1980 = {1{`RANDOM}};
  r_1995 = _RAND_1980[0:0];
  _RAND_1981 = {1{`RANDOM}};
  r_1996 = _RAND_1981[0:0];
  _RAND_1982 = {1{`RANDOM}};
  r_1997 = _RAND_1982[0:0];
  _RAND_1983 = {1{`RANDOM}};
  r_1998 = _RAND_1983[0:0];
  _RAND_1984 = {1{`RANDOM}};
  r_1999 = _RAND_1984[0:0];
  _RAND_1985 = {1{`RANDOM}};
  r_2000 = _RAND_1985[0:0];
  _RAND_1986 = {1{`RANDOM}};
  r_2001 = _RAND_1986[0:0];
  _RAND_1987 = {1{`RANDOM}};
  r_2002 = _RAND_1987[0:0];
  _RAND_1988 = {1{`RANDOM}};
  r_2003 = _RAND_1988[0:0];
  _RAND_1989 = {1{`RANDOM}};
  r_2004 = _RAND_1989[0:0];
  _RAND_1990 = {1{`RANDOM}};
  r_2005 = _RAND_1990[0:0];
  _RAND_1991 = {1{`RANDOM}};
  r_2006 = _RAND_1991[0:0];
  _RAND_1992 = {1{`RANDOM}};
  r_2007 = _RAND_1992[0:0];
  _RAND_1993 = {1{`RANDOM}};
  r_2008 = _RAND_1993[0:0];
  _RAND_1994 = {1{`RANDOM}};
  r_2009 = _RAND_1994[0:0];
  _RAND_1995 = {1{`RANDOM}};
  r_2010 = _RAND_1995[0:0];
  _RAND_1996 = {1{`RANDOM}};
  r_2011 = _RAND_1996[0:0];
  _RAND_1997 = {1{`RANDOM}};
  r_2012 = _RAND_1997[0:0];
  _RAND_1998 = {1{`RANDOM}};
  r_2013 = _RAND_1998[0:0];
  _RAND_1999 = {1{`RANDOM}};
  r_2014 = _RAND_1999[0:0];
  _RAND_2000 = {1{`RANDOM}};
  r_2015 = _RAND_2000[0:0];
  _RAND_2001 = {1{`RANDOM}};
  r_2016 = _RAND_2001[0:0];
  _RAND_2002 = {1{`RANDOM}};
  r_2017 = _RAND_2002[0:0];
  _RAND_2003 = {1{`RANDOM}};
  r_2018 = _RAND_2003[0:0];
  _RAND_2004 = {1{`RANDOM}};
  r_2019 = _RAND_2004[0:0];
  _RAND_2005 = {1{`RANDOM}};
  r_2021 = _RAND_2005[0:0];
  _RAND_2006 = {1{`RANDOM}};
  r_2022 = _RAND_2006[0:0];
  _RAND_2007 = {1{`RANDOM}};
  r_2023 = _RAND_2007[0:0];
  _RAND_2008 = {1{`RANDOM}};
  r_2024 = _RAND_2008[0:0];
  _RAND_2009 = {1{`RANDOM}};
  r_2025 = _RAND_2009[0:0];
  _RAND_2010 = {1{`RANDOM}};
  r_2026 = _RAND_2010[0:0];
  _RAND_2011 = {1{`RANDOM}};
  r_2027 = _RAND_2011[0:0];
  _RAND_2012 = {1{`RANDOM}};
  r_2028 = _RAND_2012[0:0];
  _RAND_2013 = {1{`RANDOM}};
  r_2029 = _RAND_2013[0:0];
  _RAND_2014 = {1{`RANDOM}};
  r_2030 = _RAND_2014[0:0];
  _RAND_2015 = {1{`RANDOM}};
  r_2031 = _RAND_2015[0:0];
  _RAND_2016 = {1{`RANDOM}};
  r_2032 = _RAND_2016[0:0];
  _RAND_2017 = {1{`RANDOM}};
  r_2033 = _RAND_2017[0:0];
  _RAND_2018 = {1{`RANDOM}};
  r_2034 = _RAND_2018[0:0];
  _RAND_2019 = {1{`RANDOM}};
  r_2035 = _RAND_2019[0:0];
  _RAND_2020 = {1{`RANDOM}};
  r_2036 = _RAND_2020[0:0];
  _RAND_2021 = {1{`RANDOM}};
  r_2037 = _RAND_2021[0:0];
  _RAND_2022 = {1{`RANDOM}};
  r_2038 = _RAND_2022[0:0];
  _RAND_2023 = {1{`RANDOM}};
  r_2039 = _RAND_2023[0:0];
  _RAND_2024 = {1{`RANDOM}};
  r_2040 = _RAND_2024[0:0];
  _RAND_2025 = {1{`RANDOM}};
  r_2041 = _RAND_2025[0:0];
  _RAND_2026 = {1{`RANDOM}};
  r_2042 = _RAND_2026[0:0];
  _RAND_2027 = {1{`RANDOM}};
  r_2043 = _RAND_2027[0:0];
  _RAND_2028 = {1{`RANDOM}};
  r_2044 = _RAND_2028[0:0];
  _RAND_2029 = {1{`RANDOM}};
  r_2045 = _RAND_2029[0:0];
  _RAND_2030 = {1{`RANDOM}};
  r_2046 = _RAND_2030[0:0];
  _RAND_2031 = {1{`RANDOM}};
  r_2047 = _RAND_2031[0:0];
  _RAND_2032 = {1{`RANDOM}};
  r_2048 = _RAND_2032[0:0];
  _RAND_2033 = {1{`RANDOM}};
  r_2049 = _RAND_2033[0:0];
  _RAND_2034 = {1{`RANDOM}};
  r_2050 = _RAND_2034[0:0];
  _RAND_2035 = {1{`RANDOM}};
  r_2051 = _RAND_2035[0:0];
  _RAND_2036 = {1{`RANDOM}};
  r_2052 = _RAND_2036[0:0];
  _RAND_2037 = {1{`RANDOM}};
  r_2054 = _RAND_2037[0:0];
  _RAND_2038 = {1{`RANDOM}};
  r_2055 = _RAND_2038[0:0];
  _RAND_2039 = {1{`RANDOM}};
  r_2056 = _RAND_2039[0:0];
  _RAND_2040 = {1{`RANDOM}};
  r_2057 = _RAND_2040[0:0];
  _RAND_2041 = {1{`RANDOM}};
  r_2058 = _RAND_2041[0:0];
  _RAND_2042 = {1{`RANDOM}};
  r_2059 = _RAND_2042[0:0];
  _RAND_2043 = {1{`RANDOM}};
  r_2060 = _RAND_2043[0:0];
  _RAND_2044 = {1{`RANDOM}};
  r_2061 = _RAND_2044[0:0];
  _RAND_2045 = {1{`RANDOM}};
  r_2062 = _RAND_2045[0:0];
  _RAND_2046 = {1{`RANDOM}};
  r_2063 = _RAND_2046[0:0];
  _RAND_2047 = {1{`RANDOM}};
  r_2064 = _RAND_2047[0:0];
  _RAND_2048 = {1{`RANDOM}};
  r_2065 = _RAND_2048[0:0];
  _RAND_2049 = {1{`RANDOM}};
  r_2066 = _RAND_2049[0:0];
  _RAND_2050 = {1{`RANDOM}};
  r_2067 = _RAND_2050[0:0];
  _RAND_2051 = {1{`RANDOM}};
  r_2068 = _RAND_2051[0:0];
  _RAND_2052 = {1{`RANDOM}};
  r_2069 = _RAND_2052[0:0];
  _RAND_2053 = {1{`RANDOM}};
  r_2070 = _RAND_2053[0:0];
  _RAND_2054 = {1{`RANDOM}};
  r_2071 = _RAND_2054[0:0];
  _RAND_2055 = {1{`RANDOM}};
  r_2072 = _RAND_2055[0:0];
  _RAND_2056 = {1{`RANDOM}};
  r_2073 = _RAND_2056[0:0];
  _RAND_2057 = {1{`RANDOM}};
  r_2074 = _RAND_2057[0:0];
  _RAND_2058 = {1{`RANDOM}};
  r_2075 = _RAND_2058[0:0];
  _RAND_2059 = {1{`RANDOM}};
  r_2076 = _RAND_2059[0:0];
  _RAND_2060 = {1{`RANDOM}};
  r_2077 = _RAND_2060[0:0];
  _RAND_2061 = {1{`RANDOM}};
  r_2078 = _RAND_2061[0:0];
  _RAND_2062 = {1{`RANDOM}};
  r_2079 = _RAND_2062[0:0];
  _RAND_2063 = {1{`RANDOM}};
  r_2080 = _RAND_2063[0:0];
  _RAND_2064 = {1{`RANDOM}};
  r_2081 = _RAND_2064[0:0];
  _RAND_2065 = {1{`RANDOM}};
  r_2082 = _RAND_2065[0:0];
  _RAND_2066 = {1{`RANDOM}};
  r_2083 = _RAND_2066[0:0];
  _RAND_2067 = {1{`RANDOM}};
  r_2085 = _RAND_2067[0:0];
  _RAND_2068 = {1{`RANDOM}};
  r_2086 = _RAND_2068[0:0];
  _RAND_2069 = {1{`RANDOM}};
  r_2087 = _RAND_2069[0:0];
  _RAND_2070 = {1{`RANDOM}};
  r_2088 = _RAND_2070[0:0];
  _RAND_2071 = {1{`RANDOM}};
  r_2089 = _RAND_2071[0:0];
  _RAND_2072 = {1{`RANDOM}};
  r_2090 = _RAND_2072[0:0];
  _RAND_2073 = {1{`RANDOM}};
  r_2091 = _RAND_2073[0:0];
  _RAND_2074 = {1{`RANDOM}};
  r_2092 = _RAND_2074[0:0];
  _RAND_2075 = {1{`RANDOM}};
  r_2093 = _RAND_2075[0:0];
  _RAND_2076 = {1{`RANDOM}};
  r_2094 = _RAND_2076[0:0];
  _RAND_2077 = {1{`RANDOM}};
  r_2095 = _RAND_2077[0:0];
  _RAND_2078 = {1{`RANDOM}};
  r_2096 = _RAND_2078[0:0];
  _RAND_2079 = {1{`RANDOM}};
  r_2097 = _RAND_2079[0:0];
  _RAND_2080 = {1{`RANDOM}};
  r_2098 = _RAND_2080[0:0];
  _RAND_2081 = {1{`RANDOM}};
  r_2099 = _RAND_2081[0:0];
  _RAND_2082 = {1{`RANDOM}};
  r_2100 = _RAND_2082[0:0];
  _RAND_2083 = {1{`RANDOM}};
  r_2101 = _RAND_2083[0:0];
  _RAND_2084 = {1{`RANDOM}};
  r_2102 = _RAND_2084[0:0];
  _RAND_2085 = {1{`RANDOM}};
  r_2103 = _RAND_2085[0:0];
  _RAND_2086 = {1{`RANDOM}};
  r_2104 = _RAND_2086[0:0];
  _RAND_2087 = {1{`RANDOM}};
  r_2105 = _RAND_2087[0:0];
  _RAND_2088 = {1{`RANDOM}};
  r_2106 = _RAND_2088[0:0];
  _RAND_2089 = {1{`RANDOM}};
  r_2107 = _RAND_2089[0:0];
  _RAND_2090 = {1{`RANDOM}};
  r_2108 = _RAND_2090[0:0];
  _RAND_2091 = {1{`RANDOM}};
  r_2109 = _RAND_2091[0:0];
  _RAND_2092 = {1{`RANDOM}};
  r_2110 = _RAND_2092[0:0];
  _RAND_2093 = {1{`RANDOM}};
  r_2111 = _RAND_2093[0:0];
  _RAND_2094 = {1{`RANDOM}};
  r_2112 = _RAND_2094[0:0];
  _RAND_2095 = {1{`RANDOM}};
  r_2114 = _RAND_2095[0:0];
  _RAND_2096 = {1{`RANDOM}};
  r_2115 = _RAND_2096[0:0];
  _RAND_2097 = {1{`RANDOM}};
  r_2116 = _RAND_2097[0:0];
  _RAND_2098 = {1{`RANDOM}};
  r_2117 = _RAND_2098[0:0];
  _RAND_2099 = {1{`RANDOM}};
  r_2118 = _RAND_2099[0:0];
  _RAND_2100 = {1{`RANDOM}};
  r_2119 = _RAND_2100[0:0];
  _RAND_2101 = {1{`RANDOM}};
  r_2120 = _RAND_2101[0:0];
  _RAND_2102 = {1{`RANDOM}};
  r_2121 = _RAND_2102[0:0];
  _RAND_2103 = {1{`RANDOM}};
  r_2122 = _RAND_2103[0:0];
  _RAND_2104 = {1{`RANDOM}};
  r_2123 = _RAND_2104[0:0];
  _RAND_2105 = {1{`RANDOM}};
  r_2124 = _RAND_2105[0:0];
  _RAND_2106 = {1{`RANDOM}};
  r_2125 = _RAND_2106[0:0];
  _RAND_2107 = {1{`RANDOM}};
  r_2126 = _RAND_2107[0:0];
  _RAND_2108 = {1{`RANDOM}};
  r_2127 = _RAND_2108[0:0];
  _RAND_2109 = {1{`RANDOM}};
  r_2128 = _RAND_2109[0:0];
  _RAND_2110 = {1{`RANDOM}};
  r_2129 = _RAND_2110[0:0];
  _RAND_2111 = {1{`RANDOM}};
  r_2130 = _RAND_2111[0:0];
  _RAND_2112 = {1{`RANDOM}};
  r_2131 = _RAND_2112[0:0];
  _RAND_2113 = {1{`RANDOM}};
  r_2132 = _RAND_2113[0:0];
  _RAND_2114 = {1{`RANDOM}};
  r_2133 = _RAND_2114[0:0];
  _RAND_2115 = {1{`RANDOM}};
  r_2134 = _RAND_2115[0:0];
  _RAND_2116 = {1{`RANDOM}};
  r_2135 = _RAND_2116[0:0];
  _RAND_2117 = {1{`RANDOM}};
  r_2136 = _RAND_2117[0:0];
  _RAND_2118 = {1{`RANDOM}};
  r_2137 = _RAND_2118[0:0];
  _RAND_2119 = {1{`RANDOM}};
  r_2138 = _RAND_2119[0:0];
  _RAND_2120 = {1{`RANDOM}};
  r_2139 = _RAND_2120[0:0];
  _RAND_2121 = {1{`RANDOM}};
  r_2141 = _RAND_2121[0:0];
  _RAND_2122 = {1{`RANDOM}};
  r_2142 = _RAND_2122[0:0];
  _RAND_2123 = {1{`RANDOM}};
  r_2143 = _RAND_2123[0:0];
  _RAND_2124 = {1{`RANDOM}};
  r_2144 = _RAND_2124[0:0];
  _RAND_2125 = {1{`RANDOM}};
  r_2145 = _RAND_2125[0:0];
  _RAND_2126 = {1{`RANDOM}};
  r_2146 = _RAND_2126[0:0];
  _RAND_2127 = {1{`RANDOM}};
  r_2147 = _RAND_2127[0:0];
  _RAND_2128 = {1{`RANDOM}};
  r_2148 = _RAND_2128[0:0];
  _RAND_2129 = {1{`RANDOM}};
  r_2149 = _RAND_2129[0:0];
  _RAND_2130 = {1{`RANDOM}};
  r_2150 = _RAND_2130[0:0];
  _RAND_2131 = {1{`RANDOM}};
  r_2151 = _RAND_2131[0:0];
  _RAND_2132 = {1{`RANDOM}};
  r_2152 = _RAND_2132[0:0];
  _RAND_2133 = {1{`RANDOM}};
  r_2153 = _RAND_2133[0:0];
  _RAND_2134 = {1{`RANDOM}};
  r_2154 = _RAND_2134[0:0];
  _RAND_2135 = {1{`RANDOM}};
  r_2155 = _RAND_2135[0:0];
  _RAND_2136 = {1{`RANDOM}};
  r_2156 = _RAND_2136[0:0];
  _RAND_2137 = {1{`RANDOM}};
  r_2157 = _RAND_2137[0:0];
  _RAND_2138 = {1{`RANDOM}};
  r_2158 = _RAND_2138[0:0];
  _RAND_2139 = {1{`RANDOM}};
  r_2159 = _RAND_2139[0:0];
  _RAND_2140 = {1{`RANDOM}};
  r_2160 = _RAND_2140[0:0];
  _RAND_2141 = {1{`RANDOM}};
  r_2161 = _RAND_2141[0:0];
  _RAND_2142 = {1{`RANDOM}};
  r_2162 = _RAND_2142[0:0];
  _RAND_2143 = {1{`RANDOM}};
  r_2163 = _RAND_2143[0:0];
  _RAND_2144 = {1{`RANDOM}};
  r_2164 = _RAND_2144[0:0];
  _RAND_2145 = {1{`RANDOM}};
  r_2166 = _RAND_2145[0:0];
  _RAND_2146 = {1{`RANDOM}};
  r_2167 = _RAND_2146[0:0];
  _RAND_2147 = {1{`RANDOM}};
  r_2168 = _RAND_2147[0:0];
  _RAND_2148 = {1{`RANDOM}};
  r_2169 = _RAND_2148[0:0];
  _RAND_2149 = {1{`RANDOM}};
  r_2170 = _RAND_2149[0:0];
  _RAND_2150 = {1{`RANDOM}};
  r_2171 = _RAND_2150[0:0];
  _RAND_2151 = {1{`RANDOM}};
  r_2172 = _RAND_2151[0:0];
  _RAND_2152 = {1{`RANDOM}};
  r_2173 = _RAND_2152[0:0];
  _RAND_2153 = {1{`RANDOM}};
  r_2174 = _RAND_2153[0:0];
  _RAND_2154 = {1{`RANDOM}};
  r_2175 = _RAND_2154[0:0];
  _RAND_2155 = {1{`RANDOM}};
  r_2176 = _RAND_2155[0:0];
  _RAND_2156 = {1{`RANDOM}};
  r_2177 = _RAND_2156[0:0];
  _RAND_2157 = {1{`RANDOM}};
  r_2178 = _RAND_2157[0:0];
  _RAND_2158 = {1{`RANDOM}};
  r_2179 = _RAND_2158[0:0];
  _RAND_2159 = {1{`RANDOM}};
  r_2180 = _RAND_2159[0:0];
  _RAND_2160 = {1{`RANDOM}};
  r_2181 = _RAND_2160[0:0];
  _RAND_2161 = {1{`RANDOM}};
  r_2182 = _RAND_2161[0:0];
  _RAND_2162 = {1{`RANDOM}};
  r_2183 = _RAND_2162[0:0];
  _RAND_2163 = {1{`RANDOM}};
  r_2184 = _RAND_2163[0:0];
  _RAND_2164 = {1{`RANDOM}};
  r_2185 = _RAND_2164[0:0];
  _RAND_2165 = {1{`RANDOM}};
  r_2186 = _RAND_2165[0:0];
  _RAND_2166 = {1{`RANDOM}};
  r_2187 = _RAND_2166[0:0];
  _RAND_2167 = {1{`RANDOM}};
  r_2189 = _RAND_2167[0:0];
  _RAND_2168 = {1{`RANDOM}};
  r_2190 = _RAND_2168[0:0];
  _RAND_2169 = {1{`RANDOM}};
  r_2191 = _RAND_2169[0:0];
  _RAND_2170 = {1{`RANDOM}};
  r_2192 = _RAND_2170[0:0];
  _RAND_2171 = {1{`RANDOM}};
  r_2193 = _RAND_2171[0:0];
  _RAND_2172 = {1{`RANDOM}};
  r_2194 = _RAND_2172[0:0];
  _RAND_2173 = {1{`RANDOM}};
  r_2195 = _RAND_2173[0:0];
  _RAND_2174 = {1{`RANDOM}};
  r_2196 = _RAND_2174[0:0];
  _RAND_2175 = {1{`RANDOM}};
  r_2197 = _RAND_2175[0:0];
  _RAND_2176 = {1{`RANDOM}};
  r_2198 = _RAND_2176[0:0];
  _RAND_2177 = {1{`RANDOM}};
  r_2199 = _RAND_2177[0:0];
  _RAND_2178 = {1{`RANDOM}};
  r_2200 = _RAND_2178[0:0];
  _RAND_2179 = {1{`RANDOM}};
  r_2201 = _RAND_2179[0:0];
  _RAND_2180 = {1{`RANDOM}};
  r_2202 = _RAND_2180[0:0];
  _RAND_2181 = {1{`RANDOM}};
  r_2203 = _RAND_2181[0:0];
  _RAND_2182 = {1{`RANDOM}};
  r_2204 = _RAND_2182[0:0];
  _RAND_2183 = {1{`RANDOM}};
  r_2205 = _RAND_2183[0:0];
  _RAND_2184 = {1{`RANDOM}};
  r_2206 = _RAND_2184[0:0];
  _RAND_2185 = {1{`RANDOM}};
  r_2207 = _RAND_2185[0:0];
  _RAND_2186 = {1{`RANDOM}};
  r_2208 = _RAND_2186[0:0];
  _RAND_2187 = {1{`RANDOM}};
  r_2210 = _RAND_2187[0:0];
  _RAND_2188 = {1{`RANDOM}};
  r_2211 = _RAND_2188[0:0];
  _RAND_2189 = {1{`RANDOM}};
  r_2212 = _RAND_2189[0:0];
  _RAND_2190 = {1{`RANDOM}};
  r_2213 = _RAND_2190[0:0];
  _RAND_2191 = {1{`RANDOM}};
  r_2214 = _RAND_2191[0:0];
  _RAND_2192 = {1{`RANDOM}};
  r_2215 = _RAND_2192[0:0];
  _RAND_2193 = {1{`RANDOM}};
  r_2216 = _RAND_2193[0:0];
  _RAND_2194 = {1{`RANDOM}};
  r_2217 = _RAND_2194[0:0];
  _RAND_2195 = {1{`RANDOM}};
  r_2218 = _RAND_2195[0:0];
  _RAND_2196 = {1{`RANDOM}};
  r_2219 = _RAND_2196[0:0];
  _RAND_2197 = {1{`RANDOM}};
  r_2220 = _RAND_2197[0:0];
  _RAND_2198 = {1{`RANDOM}};
  r_2221 = _RAND_2198[0:0];
  _RAND_2199 = {1{`RANDOM}};
  r_2222 = _RAND_2199[0:0];
  _RAND_2200 = {1{`RANDOM}};
  r_2223 = _RAND_2200[0:0];
  _RAND_2201 = {1{`RANDOM}};
  r_2224 = _RAND_2201[0:0];
  _RAND_2202 = {1{`RANDOM}};
  r_2225 = _RAND_2202[0:0];
  _RAND_2203 = {1{`RANDOM}};
  r_2226 = _RAND_2203[0:0];
  _RAND_2204 = {1{`RANDOM}};
  r_2227 = _RAND_2204[0:0];
  _RAND_2205 = {1{`RANDOM}};
  r_2229 = _RAND_2205[0:0];
  _RAND_2206 = {1{`RANDOM}};
  r_2230 = _RAND_2206[0:0];
  _RAND_2207 = {1{`RANDOM}};
  r_2231 = _RAND_2207[0:0];
  _RAND_2208 = {1{`RANDOM}};
  r_2232 = _RAND_2208[0:0];
  _RAND_2209 = {1{`RANDOM}};
  r_2233 = _RAND_2209[0:0];
  _RAND_2210 = {1{`RANDOM}};
  r_2234 = _RAND_2210[0:0];
  _RAND_2211 = {1{`RANDOM}};
  r_2235 = _RAND_2211[0:0];
  _RAND_2212 = {1{`RANDOM}};
  r_2236 = _RAND_2212[0:0];
  _RAND_2213 = {1{`RANDOM}};
  r_2237 = _RAND_2213[0:0];
  _RAND_2214 = {1{`RANDOM}};
  r_2238 = _RAND_2214[0:0];
  _RAND_2215 = {1{`RANDOM}};
  r_2239 = _RAND_2215[0:0];
  _RAND_2216 = {1{`RANDOM}};
  r_2240 = _RAND_2216[0:0];
  _RAND_2217 = {1{`RANDOM}};
  r_2241 = _RAND_2217[0:0];
  _RAND_2218 = {1{`RANDOM}};
  r_2242 = _RAND_2218[0:0];
  _RAND_2219 = {1{`RANDOM}};
  r_2243 = _RAND_2219[0:0];
  _RAND_2220 = {1{`RANDOM}};
  r_2244 = _RAND_2220[0:0];
  _RAND_2221 = {1{`RANDOM}};
  r_2246 = _RAND_2221[0:0];
  _RAND_2222 = {1{`RANDOM}};
  r_2247 = _RAND_2222[0:0];
  _RAND_2223 = {1{`RANDOM}};
  r_2248 = _RAND_2223[0:0];
  _RAND_2224 = {1{`RANDOM}};
  r_2249 = _RAND_2224[0:0];
  _RAND_2225 = {1{`RANDOM}};
  r_2250 = _RAND_2225[0:0];
  _RAND_2226 = {1{`RANDOM}};
  r_2251 = _RAND_2226[0:0];
  _RAND_2227 = {1{`RANDOM}};
  r_2252 = _RAND_2227[0:0];
  _RAND_2228 = {1{`RANDOM}};
  r_2253 = _RAND_2228[0:0];
  _RAND_2229 = {1{`RANDOM}};
  r_2254 = _RAND_2229[0:0];
  _RAND_2230 = {1{`RANDOM}};
  r_2255 = _RAND_2230[0:0];
  _RAND_2231 = {1{`RANDOM}};
  r_2256 = _RAND_2231[0:0];
  _RAND_2232 = {1{`RANDOM}};
  r_2257 = _RAND_2232[0:0];
  _RAND_2233 = {1{`RANDOM}};
  r_2258 = _RAND_2233[0:0];
  _RAND_2234 = {1{`RANDOM}};
  r_2259 = _RAND_2234[0:0];
  _RAND_2235 = {1{`RANDOM}};
  r_2261 = _RAND_2235[0:0];
  _RAND_2236 = {1{`RANDOM}};
  r_2262 = _RAND_2236[0:0];
  _RAND_2237 = {1{`RANDOM}};
  r_2263 = _RAND_2237[0:0];
  _RAND_2238 = {1{`RANDOM}};
  r_2264 = _RAND_2238[0:0];
  _RAND_2239 = {1{`RANDOM}};
  r_2265 = _RAND_2239[0:0];
  _RAND_2240 = {1{`RANDOM}};
  r_2266 = _RAND_2240[0:0];
  _RAND_2241 = {1{`RANDOM}};
  r_2267 = _RAND_2241[0:0];
  _RAND_2242 = {1{`RANDOM}};
  r_2268 = _RAND_2242[0:0];
  _RAND_2243 = {1{`RANDOM}};
  r_2269 = _RAND_2243[0:0];
  _RAND_2244 = {1{`RANDOM}};
  r_2270 = _RAND_2244[0:0];
  _RAND_2245 = {1{`RANDOM}};
  r_2271 = _RAND_2245[0:0];
  _RAND_2246 = {1{`RANDOM}};
  r_2272 = _RAND_2246[0:0];
  _RAND_2247 = {1{`RANDOM}};
  r_2274 = _RAND_2247[0:0];
  _RAND_2248 = {1{`RANDOM}};
  r_2275 = _RAND_2248[0:0];
  _RAND_2249 = {1{`RANDOM}};
  r_2276 = _RAND_2249[0:0];
  _RAND_2250 = {1{`RANDOM}};
  r_2277 = _RAND_2250[0:0];
  _RAND_2251 = {1{`RANDOM}};
  r_2278 = _RAND_2251[0:0];
  _RAND_2252 = {1{`RANDOM}};
  r_2279 = _RAND_2252[0:0];
  _RAND_2253 = {1{`RANDOM}};
  r_2280 = _RAND_2253[0:0];
  _RAND_2254 = {1{`RANDOM}};
  r_2281 = _RAND_2254[0:0];
  _RAND_2255 = {1{`RANDOM}};
  r_2282 = _RAND_2255[0:0];
  _RAND_2256 = {1{`RANDOM}};
  r_2283 = _RAND_2256[0:0];
  _RAND_2257 = {1{`RANDOM}};
  r_2285 = _RAND_2257[0:0];
  _RAND_2258 = {1{`RANDOM}};
  r_2286 = _RAND_2258[0:0];
  _RAND_2259 = {1{`RANDOM}};
  r_2287 = _RAND_2259[0:0];
  _RAND_2260 = {1{`RANDOM}};
  r_2288 = _RAND_2260[0:0];
  _RAND_2261 = {1{`RANDOM}};
  r_2289 = _RAND_2261[0:0];
  _RAND_2262 = {1{`RANDOM}};
  r_2290 = _RAND_2262[0:0];
  _RAND_2263 = {1{`RANDOM}};
  r_2291 = _RAND_2263[0:0];
  _RAND_2264 = {1{`RANDOM}};
  r_2292 = _RAND_2264[0:0];
  _RAND_2265 = {1{`RANDOM}};
  r_2294 = _RAND_2265[0:0];
  _RAND_2266 = {1{`RANDOM}};
  r_2295 = _RAND_2266[0:0];
  _RAND_2267 = {1{`RANDOM}};
  r_2296 = _RAND_2267[0:0];
  _RAND_2268 = {1{`RANDOM}};
  r_2297 = _RAND_2268[0:0];
  _RAND_2269 = {1{`RANDOM}};
  r_2298 = _RAND_2269[0:0];
  _RAND_2270 = {1{`RANDOM}};
  r_2299 = _RAND_2270[0:0];
  _RAND_2271 = {1{`RANDOM}};
  r_2301 = _RAND_2271[0:0];
  _RAND_2272 = {1{`RANDOM}};
  r_2302 = _RAND_2272[0:0];
  _RAND_2273 = {1{`RANDOM}};
  r_2303 = _RAND_2273[0:0];
  _RAND_2274 = {1{`RANDOM}};
  r_2304 = _RAND_2274[0:0];
  _RAND_2275 = {1{`RANDOM}};
  r_2306 = _RAND_2275[0:0];
  _RAND_2276 = {1{`RANDOM}};
  r_2307 = _RAND_2276[0:0];
  _RAND_2277 = {1{`RANDOM}};
  r_2308 = _RAND_2277[0:0];
  _RAND_2278 = {1{`RANDOM}};
  r_2309 = _RAND_2278[0:0];
  _RAND_2279 = {1{`RANDOM}};
  r_2310 = _RAND_2279[0:0];
  _RAND_2280 = {1{`RANDOM}};
  r_2311 = _RAND_2280[0:0];
  _RAND_2281 = {1{`RANDOM}};
  r_2312 = _RAND_2281[0:0];
  _RAND_2282 = {1{`RANDOM}};
  r_2313 = _RAND_2282[0:0];
  _RAND_2283 = {1{`RANDOM}};
  r_2314 = _RAND_2283[0:0];
  _RAND_2284 = {1{`RANDOM}};
  r_2315 = _RAND_2284[0:0];
  _RAND_2285 = {1{`RANDOM}};
  r_2316 = _RAND_2285[0:0];
  _RAND_2286 = {1{`RANDOM}};
  r_2317 = _RAND_2286[0:0];
  _RAND_2287 = {1{`RANDOM}};
  r_2318 = _RAND_2287[0:0];
  _RAND_2288 = {1{`RANDOM}};
  r_2319 = _RAND_2288[0:0];
  _RAND_2289 = {1{`RANDOM}};
  r_2320 = _RAND_2289[0:0];
  _RAND_2290 = {1{`RANDOM}};
  r_2321 = _RAND_2290[0:0];
  _RAND_2291 = {1{`RANDOM}};
  r_2322 = _RAND_2291[0:0];
  _RAND_2292 = {1{`RANDOM}};
  r_2323 = _RAND_2292[0:0];
  _RAND_2293 = {1{`RANDOM}};
  r_2324 = _RAND_2293[0:0];
  _RAND_2294 = {1{`RANDOM}};
  r_2325 = _RAND_2294[0:0];
  _RAND_2295 = {1{`RANDOM}};
  r_2326 = _RAND_2295[0:0];
  _RAND_2296 = {1{`RANDOM}};
  r_2327 = _RAND_2296[0:0];
  _RAND_2297 = {1{`RANDOM}};
  r_2328 = _RAND_2297[0:0];
  _RAND_2298 = {1{`RANDOM}};
  r_2329 = _RAND_2298[0:0];
  _RAND_2299 = {1{`RANDOM}};
  r_2330 = _RAND_2299[0:0];
  _RAND_2300 = {1{`RANDOM}};
  r_2331 = _RAND_2300[0:0];
  _RAND_2301 = {1{`RANDOM}};
  r_2332 = _RAND_2301[0:0];
  _RAND_2302 = {1{`RANDOM}};
  r_2333 = _RAND_2302[0:0];
  _RAND_2303 = {1{`RANDOM}};
  r_2334 = _RAND_2303[0:0];
  _RAND_2304 = {1{`RANDOM}};
  r_2335 = _RAND_2304[0:0];
  _RAND_2305 = {1{`RANDOM}};
  r_2336 = _RAND_2305[0:0];
  _RAND_2306 = {1{`RANDOM}};
  r_2337 = _RAND_2306[0:0];
  _RAND_2307 = {1{`RANDOM}};
  r_2338 = _RAND_2307[0:0];
  _RAND_2308 = {1{`RANDOM}};
  r_2339 = _RAND_2308[0:0];
  _RAND_2309 = {1{`RANDOM}};
  r_2340 = _RAND_2309[0:0];
  _RAND_2310 = {1{`RANDOM}};
  r_2341 = _RAND_2310[0:0];
  _RAND_2311 = {1{`RANDOM}};
  r_2342 = _RAND_2311[0:0];
  _RAND_2312 = {1{`RANDOM}};
  r_2343 = _RAND_2312[0:0];
  _RAND_2313 = {1{`RANDOM}};
  r_2344 = _RAND_2313[0:0];
  _RAND_2314 = {1{`RANDOM}};
  r_2345 = _RAND_2314[0:0];
  _RAND_2315 = {1{`RANDOM}};
  r_2346 = _RAND_2315[0:0];
  _RAND_2316 = {1{`RANDOM}};
  r_2347 = _RAND_2316[0:0];
  _RAND_2317 = {1{`RANDOM}};
  r_2348 = _RAND_2317[0:0];
  _RAND_2318 = {1{`RANDOM}};
  r_2349 = _RAND_2318[0:0];
  _RAND_2319 = {1{`RANDOM}};
  r_2350 = _RAND_2319[0:0];
  _RAND_2320 = {1{`RANDOM}};
  r_2351 = _RAND_2320[0:0];
  _RAND_2321 = {1{`RANDOM}};
  r_2352 = _RAND_2321[0:0];
  _RAND_2322 = {1{`RANDOM}};
  r_2353 = _RAND_2322[0:0];
  _RAND_2323 = {1{`RANDOM}};
  r_2354 = _RAND_2323[0:0];
  _RAND_2324 = {1{`RANDOM}};
  r_2355 = _RAND_2324[0:0];
  _RAND_2325 = {1{`RANDOM}};
  r_2356 = _RAND_2325[0:0];
  _RAND_2326 = {1{`RANDOM}};
  r_2357 = _RAND_2326[0:0];
  _RAND_2327 = {1{`RANDOM}};
  r_2358 = _RAND_2327[0:0];
  _RAND_2328 = {1{`RANDOM}};
  r_2359 = _RAND_2328[0:0];
  _RAND_2329 = {1{`RANDOM}};
  r_2360 = _RAND_2329[0:0];
  _RAND_2330 = {1{`RANDOM}};
  r_2361 = _RAND_2330[0:0];
  _RAND_2331 = {1{`RANDOM}};
  r_2362 = _RAND_2331[0:0];
  _RAND_2332 = {1{`RANDOM}};
  r_2363 = _RAND_2332[0:0];
  _RAND_2333 = {1{`RANDOM}};
  r_2364 = _RAND_2333[0:0];
  _RAND_2334 = {1{`RANDOM}};
  r_2365 = _RAND_2334[0:0];
  _RAND_2335 = {1{`RANDOM}};
  r_2366 = _RAND_2335[0:0];
  _RAND_2336 = {1{`RANDOM}};
  r_2367 = _RAND_2336[0:0];
  _RAND_2337 = {1{`RANDOM}};
  r_2368 = _RAND_2337[0:0];
  _RAND_2338 = {1{`RANDOM}};
  r_2369 = _RAND_2338[0:0];
  _RAND_2339 = {1{`RANDOM}};
  r_2370 = _RAND_2339[0:0];
  _RAND_2340 = {1{`RANDOM}};
  r_2371 = _RAND_2340[0:0];
  _RAND_2341 = {1{`RANDOM}};
  r_2372 = _RAND_2341[0:0];
  _RAND_2342 = {1{`RANDOM}};
  r_2373 = _RAND_2342[0:0];
  _RAND_2343 = {1{`RANDOM}};
  r_2374 = _RAND_2343[0:0];
  _RAND_2344 = {1{`RANDOM}};
  r_2375 = _RAND_2344[0:0];
  _RAND_2345 = {1{`RANDOM}};
  r_2376 = _RAND_2345[0:0];
  _RAND_2346 = {1{`RANDOM}};
  r_2377 = _RAND_2346[0:0];
  _RAND_2347 = {1{`RANDOM}};
  r_2378 = _RAND_2347[0:0];
  _RAND_2348 = {1{`RANDOM}};
  r_2379 = _RAND_2348[0:0];
  _RAND_2349 = {1{`RANDOM}};
  r_2380 = _RAND_2349[0:0];
  _RAND_2350 = {1{`RANDOM}};
  r_2381 = _RAND_2350[0:0];
  _RAND_2351 = {1{`RANDOM}};
  r_2382 = _RAND_2351[0:0];
  _RAND_2352 = {1{`RANDOM}};
  r_2383 = _RAND_2352[0:0];
  _RAND_2353 = {1{`RANDOM}};
  r_2384 = _RAND_2353[0:0];
  _RAND_2354 = {1{`RANDOM}};
  r_2385 = _RAND_2354[0:0];
  _RAND_2355 = {1{`RANDOM}};
  r_2386 = _RAND_2355[0:0];
  _RAND_2356 = {1{`RANDOM}};
  r_2387 = _RAND_2356[0:0];
  _RAND_2357 = {1{`RANDOM}};
  r_2388 = _RAND_2357[0:0];
  _RAND_2358 = {1{`RANDOM}};
  r_2389 = _RAND_2358[0:0];
  _RAND_2359 = {1{`RANDOM}};
  r_2390 = _RAND_2359[0:0];
  _RAND_2360 = {1{`RANDOM}};
  r_2391 = _RAND_2360[0:0];
  _RAND_2361 = {1{`RANDOM}};
  r_2392 = _RAND_2361[0:0];
  _RAND_2362 = {1{`RANDOM}};
  r_2393 = _RAND_2362[0:0];
  _RAND_2363 = {1{`RANDOM}};
  r_2394 = _RAND_2363[0:0];
  _RAND_2364 = {1{`RANDOM}};
  r_2395 = _RAND_2364[0:0];
  _RAND_2365 = {1{`RANDOM}};
  r_2396 = _RAND_2365[0:0];
  _RAND_2366 = {1{`RANDOM}};
  r_2397 = _RAND_2366[0:0];
  _RAND_2367 = {1{`RANDOM}};
  r_2398 = _RAND_2367[0:0];
  _RAND_2368 = {1{`RANDOM}};
  r_2399 = _RAND_2368[0:0];
  _RAND_2369 = {1{`RANDOM}};
  r_2400 = _RAND_2369[0:0];
  _RAND_2370 = {1{`RANDOM}};
  r_2401 = _RAND_2370[0:0];
  _RAND_2371 = {1{`RANDOM}};
  r_2402 = _RAND_2371[0:0];
  _RAND_2372 = {1{`RANDOM}};
  r_2403 = _RAND_2372[0:0];
  _RAND_2373 = {1{`RANDOM}};
  r_2404 = _RAND_2373[0:0];
  _RAND_2374 = {1{`RANDOM}};
  r_2405 = _RAND_2374[0:0];
  _RAND_2375 = {1{`RANDOM}};
  r_2406 = _RAND_2375[0:0];
  _RAND_2376 = {1{`RANDOM}};
  r_2407 = _RAND_2376[0:0];
  _RAND_2377 = {1{`RANDOM}};
  r_2408 = _RAND_2377[0:0];
  _RAND_2378 = {1{`RANDOM}};
  r_2409 = _RAND_2378[0:0];
  _RAND_2379 = {1{`RANDOM}};
  r_2410 = _RAND_2379[0:0];
  _RAND_2380 = {1{`RANDOM}};
  r_2411 = _RAND_2380[0:0];
  _RAND_2381 = {1{`RANDOM}};
  r_2412 = _RAND_2381[0:0];
  _RAND_2382 = {1{`RANDOM}};
  r_2413 = _RAND_2382[0:0];
  _RAND_2383 = {1{`RANDOM}};
  r_2414 = _RAND_2383[0:0];
  _RAND_2384 = {1{`RANDOM}};
  r_2415 = _RAND_2384[0:0];
  _RAND_2385 = {1{`RANDOM}};
  r_2416 = _RAND_2385[0:0];
  _RAND_2386 = {1{`RANDOM}};
  r_2417 = _RAND_2386[0:0];
  _RAND_2387 = {1{`RANDOM}};
  r_2418 = _RAND_2387[0:0];
  _RAND_2388 = {1{`RANDOM}};
  r_2419 = _RAND_2388[0:0];
  _RAND_2389 = {1{`RANDOM}};
  r_2420 = _RAND_2389[0:0];
  _RAND_2390 = {1{`RANDOM}};
  r_2421 = _RAND_2390[0:0];
  _RAND_2391 = {1{`RANDOM}};
  r_2422 = _RAND_2391[0:0];
  _RAND_2392 = {1{`RANDOM}};
  r_2423 = _RAND_2392[0:0];
  _RAND_2393 = {1{`RANDOM}};
  r_2424 = _RAND_2393[0:0];
  _RAND_2394 = {1{`RANDOM}};
  r_2425 = _RAND_2394[0:0];
  _RAND_2395 = {1{`RANDOM}};
  r_2426 = _RAND_2395[0:0];
  _RAND_2396 = {1{`RANDOM}};
  r_2427 = _RAND_2396[0:0];
  _RAND_2397 = {1{`RANDOM}};
  r_2428 = _RAND_2397[0:0];
  _RAND_2398 = {1{`RANDOM}};
  r_2429 = _RAND_2398[0:0];
  _RAND_2399 = {1{`RANDOM}};
  r_2430 = _RAND_2399[0:0];
  _RAND_2400 = {1{`RANDOM}};
  r_2431 = _RAND_2400[0:0];
  _RAND_2401 = {1{`RANDOM}};
  r_2432 = _RAND_2401[0:0];
  _RAND_2402 = {1{`RANDOM}};
  r_2433 = _RAND_2402[0:0];
  _RAND_2403 = {1{`RANDOM}};
  r_2434 = _RAND_2403[0:0];
  _RAND_2404 = {1{`RANDOM}};
  r_2435 = _RAND_2404[0:0];
  _RAND_2405 = {1{`RANDOM}};
  r_2436 = _RAND_2405[0:0];
  _RAND_2406 = {1{`RANDOM}};
  r_2437 = _RAND_2406[0:0];
  _RAND_2407 = {1{`RANDOM}};
  r_2438 = _RAND_2407[0:0];
  _RAND_2408 = {1{`RANDOM}};
  r_2439 = _RAND_2408[0:0];
  _RAND_2409 = {1{`RANDOM}};
  r_2440 = _RAND_2409[0:0];
  _RAND_2410 = {1{`RANDOM}};
  r_2441 = _RAND_2410[0:0];
  _RAND_2411 = {1{`RANDOM}};
  r_2442 = _RAND_2411[0:0];
  _RAND_2412 = {1{`RANDOM}};
  r_2443 = _RAND_2412[0:0];
  _RAND_2413 = {1{`RANDOM}};
  r_2444 = _RAND_2413[0:0];
  _RAND_2414 = {1{`RANDOM}};
  r_2445 = _RAND_2414[0:0];
  _RAND_2415 = {1{`RANDOM}};
  r_2446 = _RAND_2415[0:0];
  _RAND_2416 = {1{`RANDOM}};
  r_2447 = _RAND_2416[0:0];
  _RAND_2417 = {1{`RANDOM}};
  r_2448 = _RAND_2417[0:0];
  _RAND_2418 = {1{`RANDOM}};
  r_2449 = _RAND_2418[0:0];
  _RAND_2419 = {1{`RANDOM}};
  r_2450 = _RAND_2419[0:0];
  _RAND_2420 = {1{`RANDOM}};
  r_2451 = _RAND_2420[0:0];
  _RAND_2421 = {1{`RANDOM}};
  r_2452 = _RAND_2421[0:0];
  _RAND_2422 = {1{`RANDOM}};
  r_2453 = _RAND_2422[0:0];
  _RAND_2423 = {1{`RANDOM}};
  r_2454 = _RAND_2423[0:0];
  _RAND_2424 = {1{`RANDOM}};
  r_2455 = _RAND_2424[0:0];
  _RAND_2425 = {1{`RANDOM}};
  r_2456 = _RAND_2425[0:0];
  _RAND_2426 = {1{`RANDOM}};
  r_2457 = _RAND_2426[0:0];
  _RAND_2427 = {1{`RANDOM}};
  r_2458 = _RAND_2427[0:0];
  _RAND_2428 = {1{`RANDOM}};
  r_2459 = _RAND_2428[0:0];
  _RAND_2429 = {1{`RANDOM}};
  r_2460 = _RAND_2429[0:0];
  _RAND_2430 = {1{`RANDOM}};
  r_2461 = _RAND_2430[0:0];
  _RAND_2431 = {1{`RANDOM}};
  r_2462 = _RAND_2431[0:0];
  _RAND_2432 = {1{`RANDOM}};
  r_2463 = _RAND_2432[0:0];
  _RAND_2433 = {1{`RANDOM}};
  r_2464 = _RAND_2433[0:0];
  _RAND_2434 = {1{`RANDOM}};
  r_2465 = _RAND_2434[0:0];
  _RAND_2435 = {1{`RANDOM}};
  r_2466 = _RAND_2435[0:0];
  _RAND_2436 = {1{`RANDOM}};
  r_2467 = _RAND_2436[0:0];
  _RAND_2437 = {1{`RANDOM}};
  r_2468 = _RAND_2437[0:0];
  _RAND_2438 = {1{`RANDOM}};
  r_2469 = _RAND_2438[0:0];
  _RAND_2439 = {1{`RANDOM}};
  r_2470 = _RAND_2439[0:0];
  _RAND_2440 = {1{`RANDOM}};
  r_2471 = _RAND_2440[0:0];
  _RAND_2441 = {1{`RANDOM}};
  r_2472 = _RAND_2441[0:0];
  _RAND_2442 = {1{`RANDOM}};
  r_2473 = _RAND_2442[0:0];
  _RAND_2443 = {1{`RANDOM}};
  r_2474 = _RAND_2443[0:0];
  _RAND_2444 = {1{`RANDOM}};
  r_2475 = _RAND_2444[0:0];
  _RAND_2445 = {1{`RANDOM}};
  r_2476 = _RAND_2445[0:0];
  _RAND_2446 = {1{`RANDOM}};
  r_2477 = _RAND_2446[0:0];
  _RAND_2447 = {1{`RANDOM}};
  r_2478 = _RAND_2447[0:0];
  _RAND_2448 = {1{`RANDOM}};
  r_2479 = _RAND_2448[0:0];
  _RAND_2449 = {1{`RANDOM}};
  r_2480 = _RAND_2449[0:0];
  _RAND_2450 = {1{`RANDOM}};
  r_2481 = _RAND_2450[0:0];
  _RAND_2451 = {1{`RANDOM}};
  r_2482 = _RAND_2451[0:0];
  _RAND_2452 = {1{`RANDOM}};
  r_2483 = _RAND_2452[0:0];
  _RAND_2453 = {1{`RANDOM}};
  r_2484 = _RAND_2453[0:0];
  _RAND_2454 = {1{`RANDOM}};
  r_2485 = _RAND_2454[0:0];
  _RAND_2455 = {1{`RANDOM}};
  r_2486 = _RAND_2455[0:0];
  _RAND_2456 = {1{`RANDOM}};
  r_2487 = _RAND_2456[0:0];
  _RAND_2457 = {1{`RANDOM}};
  r_2488 = _RAND_2457[0:0];
  _RAND_2458 = {1{`RANDOM}};
  r_2489 = _RAND_2458[0:0];
  _RAND_2459 = {1{`RANDOM}};
  r_2490 = _RAND_2459[0:0];
  _RAND_2460 = {1{`RANDOM}};
  r_2491 = _RAND_2460[0:0];
  _RAND_2461 = {1{`RANDOM}};
  r_2492 = _RAND_2461[0:0];
  _RAND_2462 = {1{`RANDOM}};
  r_2493 = _RAND_2462[0:0];
  _RAND_2463 = {1{`RANDOM}};
  r_2494 = _RAND_2463[0:0];
  _RAND_2464 = {1{`RANDOM}};
  r_2495 = _RAND_2464[0:0];
  _RAND_2465 = {1{`RANDOM}};
  r_2496 = _RAND_2465[0:0];
  _RAND_2466 = {1{`RANDOM}};
  r_2497 = _RAND_2466[0:0];
  _RAND_2467 = {1{`RANDOM}};
  r_2498 = _RAND_2467[0:0];
  _RAND_2468 = {1{`RANDOM}};
  r_2499 = _RAND_2468[0:0];
  _RAND_2469 = {1{`RANDOM}};
  r_2500 = _RAND_2469[0:0];
  _RAND_2470 = {1{`RANDOM}};
  r_2501 = _RAND_2470[0:0];
  _RAND_2471 = {1{`RANDOM}};
  r_2502 = _RAND_2471[0:0];
  _RAND_2472 = {1{`RANDOM}};
  r_2503 = _RAND_2472[0:0];
  _RAND_2473 = {1{`RANDOM}};
  r_2504 = _RAND_2473[0:0];
  _RAND_2474 = {1{`RANDOM}};
  r_2505 = _RAND_2474[0:0];
  _RAND_2475 = {1{`RANDOM}};
  r_2506 = _RAND_2475[0:0];
  _RAND_2476 = {1{`RANDOM}};
  r_2507 = _RAND_2476[0:0];
  _RAND_2477 = {1{`RANDOM}};
  r_2508 = _RAND_2477[0:0];
  _RAND_2478 = {1{`RANDOM}};
  r_2509 = _RAND_2478[0:0];
  _RAND_2479 = {1{`RANDOM}};
  r_2510 = _RAND_2479[0:0];
  _RAND_2480 = {1{`RANDOM}};
  r_2511 = _RAND_2480[0:0];
  _RAND_2481 = {1{`RANDOM}};
  r_2512 = _RAND_2481[0:0];
  _RAND_2482 = {1{`RANDOM}};
  r_2513 = _RAND_2482[0:0];
  _RAND_2483 = {1{`RANDOM}};
  r_2514 = _RAND_2483[0:0];
  _RAND_2484 = {1{`RANDOM}};
  r_2515 = _RAND_2484[0:0];
  _RAND_2485 = {1{`RANDOM}};
  r_2516 = _RAND_2485[0:0];
  _RAND_2486 = {1{`RANDOM}};
  r_2517 = _RAND_2486[0:0];
  _RAND_2487 = {1{`RANDOM}};
  r_2518 = _RAND_2487[0:0];
  _RAND_2488 = {1{`RANDOM}};
  r_2519 = _RAND_2488[0:0];
  _RAND_2489 = {1{`RANDOM}};
  r_2520 = _RAND_2489[0:0];
  _RAND_2490 = {1{`RANDOM}};
  r_2521 = _RAND_2490[0:0];
  _RAND_2491 = {1{`RANDOM}};
  r_2522 = _RAND_2491[0:0];
  _RAND_2492 = {1{`RANDOM}};
  r_2523 = _RAND_2492[0:0];
  _RAND_2493 = {1{`RANDOM}};
  r_2524 = _RAND_2493[0:0];
  _RAND_2494 = {1{`RANDOM}};
  r_2525 = _RAND_2494[0:0];
  _RAND_2495 = {1{`RANDOM}};
  r_2526 = _RAND_2495[0:0];
  _RAND_2496 = {1{`RANDOM}};
  r_2527 = _RAND_2496[0:0];
  _RAND_2497 = {1{`RANDOM}};
  r_2528 = _RAND_2497[0:0];
  _RAND_2498 = {1{`RANDOM}};
  r_2529 = _RAND_2498[0:0];
  _RAND_2499 = {1{`RANDOM}};
  r_2530 = _RAND_2499[0:0];
  _RAND_2500 = {1{`RANDOM}};
  r_2531 = _RAND_2500[0:0];
  _RAND_2501 = {1{`RANDOM}};
  r_2532 = _RAND_2501[0:0];
  _RAND_2502 = {1{`RANDOM}};
  r_2533 = _RAND_2502[0:0];
  _RAND_2503 = {1{`RANDOM}};
  r_2534 = _RAND_2503[0:0];
  _RAND_2504 = {1{`RANDOM}};
  r_2535 = _RAND_2504[0:0];
  _RAND_2505 = {1{`RANDOM}};
  r_2536 = _RAND_2505[0:0];
  _RAND_2506 = {1{`RANDOM}};
  r_2537 = _RAND_2506[0:0];
  _RAND_2507 = {1{`RANDOM}};
  r_2538 = _RAND_2507[0:0];
  _RAND_2508 = {1{`RANDOM}};
  r_2539 = _RAND_2508[0:0];
  _RAND_2509 = {1{`RANDOM}};
  r_2540 = _RAND_2509[0:0];
  _RAND_2510 = {1{`RANDOM}};
  r_2541 = _RAND_2510[0:0];
  _RAND_2511 = {1{`RANDOM}};
  r_2542 = _RAND_2511[0:0];
  _RAND_2512 = {1{`RANDOM}};
  r_2543 = _RAND_2512[0:0];
  _RAND_2513 = {1{`RANDOM}};
  r_2544 = _RAND_2513[0:0];
  _RAND_2514 = {1{`RANDOM}};
  r_2545 = _RAND_2514[0:0];
  _RAND_2515 = {1{`RANDOM}};
  r_2546 = _RAND_2515[0:0];
  _RAND_2516 = {1{`RANDOM}};
  r_2547 = _RAND_2516[0:0];
  _RAND_2517 = {1{`RANDOM}};
  r_2548 = _RAND_2517[0:0];
  _RAND_2518 = {1{`RANDOM}};
  r_2549 = _RAND_2518[0:0];
  _RAND_2519 = {1{`RANDOM}};
  r_2550 = _RAND_2519[0:0];
  _RAND_2520 = {1{`RANDOM}};
  r_2551 = _RAND_2520[0:0];
  _RAND_2521 = {1{`RANDOM}};
  r_2552 = _RAND_2521[0:0];
  _RAND_2522 = {1{`RANDOM}};
  r_2553 = _RAND_2522[0:0];
  _RAND_2523 = {1{`RANDOM}};
  r_2554 = _RAND_2523[0:0];
  _RAND_2524 = {1{`RANDOM}};
  r_2555 = _RAND_2524[0:0];
  _RAND_2525 = {1{`RANDOM}};
  r_2556 = _RAND_2525[0:0];
  _RAND_2526 = {1{`RANDOM}};
  r_2557 = _RAND_2526[0:0];
  _RAND_2527 = {1{`RANDOM}};
  r_2558 = _RAND_2527[0:0];
  _RAND_2528 = {1{`RANDOM}};
  r_2559 = _RAND_2528[0:0];
  _RAND_2529 = {1{`RANDOM}};
  r_2560 = _RAND_2529[0:0];
  _RAND_2530 = {1{`RANDOM}};
  r_2561 = _RAND_2530[0:0];
  _RAND_2531 = {1{`RANDOM}};
  r_2562 = _RAND_2531[0:0];
  _RAND_2532 = {1{`RANDOM}};
  r_2563 = _RAND_2532[0:0];
  _RAND_2533 = {1{`RANDOM}};
  r_2564 = _RAND_2533[0:0];
  _RAND_2534 = {1{`RANDOM}};
  r_2565 = _RAND_2534[0:0];
  _RAND_2535 = {1{`RANDOM}};
  r_2566 = _RAND_2535[0:0];
  _RAND_2536 = {1{`RANDOM}};
  r_2567 = _RAND_2536[0:0];
  _RAND_2537 = {1{`RANDOM}};
  r_2568 = _RAND_2537[0:0];
  _RAND_2538 = {1{`RANDOM}};
  r_2569 = _RAND_2538[0:0];
  _RAND_2539 = {1{`RANDOM}};
  r_2570 = _RAND_2539[0:0];
  _RAND_2540 = {1{`RANDOM}};
  r_2571 = _RAND_2540[0:0];
  _RAND_2541 = {1{`RANDOM}};
  r_2572 = _RAND_2541[0:0];
  _RAND_2542 = {1{`RANDOM}};
  r_2573 = _RAND_2542[0:0];
  _RAND_2543 = {1{`RANDOM}};
  r_2574 = _RAND_2543[0:0];
  _RAND_2544 = {1{`RANDOM}};
  r_2575 = _RAND_2544[0:0];
  _RAND_2545 = {1{`RANDOM}};
  r_2576 = _RAND_2545[0:0];
  _RAND_2546 = {1{`RANDOM}};
  r_2577 = _RAND_2546[0:0];
  _RAND_2547 = {1{`RANDOM}};
  r_2578 = _RAND_2547[0:0];
  _RAND_2548 = {1{`RANDOM}};
  r_2579 = _RAND_2548[0:0];
  _RAND_2549 = {1{`RANDOM}};
  r_2580 = _RAND_2549[0:0];
  _RAND_2550 = {1{`RANDOM}};
  r_2581 = _RAND_2550[0:0];
  _RAND_2551 = {1{`RANDOM}};
  r_2582 = _RAND_2551[0:0];
  _RAND_2552 = {1{`RANDOM}};
  r_2583 = _RAND_2552[0:0];
  _RAND_2553 = {1{`RANDOM}};
  r_2584 = _RAND_2553[0:0];
  _RAND_2554 = {1{`RANDOM}};
  r_2585 = _RAND_2554[0:0];
  _RAND_2555 = {1{`RANDOM}};
  r_2586 = _RAND_2555[0:0];
  _RAND_2556 = {1{`RANDOM}};
  r_2587 = _RAND_2556[0:0];
  _RAND_2557 = {1{`RANDOM}};
  r_2588 = _RAND_2557[0:0];
  _RAND_2558 = {1{`RANDOM}};
  r_2589 = _RAND_2558[0:0];
  _RAND_2559 = {1{`RANDOM}};
  r_2590 = _RAND_2559[0:0];
  _RAND_2560 = {1{`RANDOM}};
  r_2591 = _RAND_2560[0:0];
  _RAND_2561 = {1{`RANDOM}};
  r_2592 = _RAND_2561[0:0];
  _RAND_2562 = {1{`RANDOM}};
  r_2593 = _RAND_2562[0:0];
  _RAND_2563 = {1{`RANDOM}};
  r_2594 = _RAND_2563[0:0];
  _RAND_2564 = {1{`RANDOM}};
  r_2595 = _RAND_2564[0:0];
  _RAND_2565 = {1{`RANDOM}};
  r_2596 = _RAND_2565[0:0];
  _RAND_2566 = {1{`RANDOM}};
  r_2597 = _RAND_2566[0:0];
  _RAND_2567 = {1{`RANDOM}};
  r_2598 = _RAND_2567[0:0];
  _RAND_2568 = {1{`RANDOM}};
  r_2599 = _RAND_2568[0:0];
  _RAND_2569 = {1{`RANDOM}};
  r_2600 = _RAND_2569[0:0];
  _RAND_2570 = {1{`RANDOM}};
  r_2601 = _RAND_2570[0:0];
  _RAND_2571 = {1{`RANDOM}};
  r_2602 = _RAND_2571[0:0];
  _RAND_2572 = {1{`RANDOM}};
  r_2603 = _RAND_2572[0:0];
  _RAND_2573 = {1{`RANDOM}};
  r_2604 = _RAND_2573[0:0];
  _RAND_2574 = {1{`RANDOM}};
  r_2605 = _RAND_2574[0:0];
  _RAND_2575 = {1{`RANDOM}};
  r_2606 = _RAND_2575[0:0];
  _RAND_2576 = {1{`RANDOM}};
  r_2607 = _RAND_2576[0:0];
  _RAND_2577 = {1{`RANDOM}};
  r_2608 = _RAND_2577[0:0];
  _RAND_2578 = {1{`RANDOM}};
  r_2609 = _RAND_2578[0:0];
  _RAND_2579 = {1{`RANDOM}};
  r_2610 = _RAND_2579[0:0];
  _RAND_2580 = {1{`RANDOM}};
  r_2611 = _RAND_2580[0:0];
  _RAND_2581 = {1{`RANDOM}};
  r_2612 = _RAND_2581[0:0];
  _RAND_2582 = {1{`RANDOM}};
  r_2613 = _RAND_2582[0:0];
  _RAND_2583 = {1{`RANDOM}};
  r_2614 = _RAND_2583[0:0];
  _RAND_2584 = {1{`RANDOM}};
  r_2615 = _RAND_2584[0:0];
  _RAND_2585 = {1{`RANDOM}};
  r_2616 = _RAND_2585[0:0];
  _RAND_2586 = {1{`RANDOM}};
  r_2617 = _RAND_2586[0:0];
  _RAND_2587 = {1{`RANDOM}};
  r_2618 = _RAND_2587[0:0];
  _RAND_2588 = {1{`RANDOM}};
  r_2619 = _RAND_2588[0:0];
  _RAND_2589 = {1{`RANDOM}};
  r_2620 = _RAND_2589[0:0];
  _RAND_2590 = {1{`RANDOM}};
  r_2621 = _RAND_2590[0:0];
  _RAND_2591 = {1{`RANDOM}};
  r_2622 = _RAND_2591[0:0];
  _RAND_2592 = {1{`RANDOM}};
  r_2623 = _RAND_2592[0:0];
  _RAND_2593 = {1{`RANDOM}};
  r_2624 = _RAND_2593[0:0];
  _RAND_2594 = {1{`RANDOM}};
  r_2625 = _RAND_2594[0:0];
  _RAND_2595 = {1{`RANDOM}};
  r_2626 = _RAND_2595[0:0];
  _RAND_2596 = {1{`RANDOM}};
  r_2627 = _RAND_2596[0:0];
  _RAND_2597 = {1{`RANDOM}};
  r_2628 = _RAND_2597[0:0];
  _RAND_2598 = {1{`RANDOM}};
  r_2629 = _RAND_2598[0:0];
  _RAND_2599 = {1{`RANDOM}};
  r_2630 = _RAND_2599[0:0];
  _RAND_2600 = {1{`RANDOM}};
  r_2631 = _RAND_2600[0:0];
  _RAND_2601 = {1{`RANDOM}};
  r_2632 = _RAND_2601[0:0];
  _RAND_2602 = {1{`RANDOM}};
  r_2633 = _RAND_2602[0:0];
  _RAND_2603 = {1{`RANDOM}};
  r_2634 = _RAND_2603[0:0];
  _RAND_2604 = {1{`RANDOM}};
  r_2635 = _RAND_2604[0:0];
  _RAND_2605 = {1{`RANDOM}};
  r_2636 = _RAND_2605[0:0];
  _RAND_2606 = {1{`RANDOM}};
  r_2637 = _RAND_2606[0:0];
  _RAND_2607 = {1{`RANDOM}};
  r_2638 = _RAND_2607[0:0];
  _RAND_2608 = {1{`RANDOM}};
  r_2639 = _RAND_2608[0:0];
  _RAND_2609 = {1{`RANDOM}};
  r_2640 = _RAND_2609[0:0];
  _RAND_2610 = {1{`RANDOM}};
  r_2641 = _RAND_2610[0:0];
  _RAND_2611 = {1{`RANDOM}};
  r_2642 = _RAND_2611[0:0];
  _RAND_2612 = {1{`RANDOM}};
  r_2643 = _RAND_2612[0:0];
  _RAND_2613 = {1{`RANDOM}};
  r_2644 = _RAND_2613[0:0];
  _RAND_2614 = {1{`RANDOM}};
  r_2645 = _RAND_2614[0:0];
  _RAND_2615 = {1{`RANDOM}};
  r_2646 = _RAND_2615[0:0];
  _RAND_2616 = {1{`RANDOM}};
  r_2647 = _RAND_2616[0:0];
  _RAND_2617 = {1{`RANDOM}};
  r_2648 = _RAND_2617[0:0];
  _RAND_2618 = {1{`RANDOM}};
  r_2649 = _RAND_2618[0:0];
  _RAND_2619 = {1{`RANDOM}};
  r_2650 = _RAND_2619[0:0];
  _RAND_2620 = {1{`RANDOM}};
  r_2651 = _RAND_2620[0:0];
  _RAND_2621 = {1{`RANDOM}};
  r_2652 = _RAND_2621[0:0];
  _RAND_2622 = {1{`RANDOM}};
  r_2653 = _RAND_2622[0:0];
  _RAND_2623 = {1{`RANDOM}};
  r_2654 = _RAND_2623[0:0];
  _RAND_2624 = {1{`RANDOM}};
  r_2655 = _RAND_2624[0:0];
  _RAND_2625 = {1{`RANDOM}};
  r_2656 = _RAND_2625[0:0];
  _RAND_2626 = {1{`RANDOM}};
  r_2657 = _RAND_2626[0:0];
  _RAND_2627 = {1{`RANDOM}};
  r_2658 = _RAND_2627[0:0];
  _RAND_2628 = {1{`RANDOM}};
  r_2659 = _RAND_2628[0:0];
  _RAND_2629 = {1{`RANDOM}};
  r_2660 = _RAND_2629[0:0];
  _RAND_2630 = {1{`RANDOM}};
  r_2661 = _RAND_2630[0:0];
  _RAND_2631 = {1{`RANDOM}};
  r_2662 = _RAND_2631[0:0];
  _RAND_2632 = {1{`RANDOM}};
  r_2663 = _RAND_2632[0:0];
  _RAND_2633 = {1{`RANDOM}};
  r_2664 = _RAND_2633[0:0];
  _RAND_2634 = {1{`RANDOM}};
  r_2665 = _RAND_2634[0:0];
  _RAND_2635 = {1{`RANDOM}};
  r_2666 = _RAND_2635[0:0];
  _RAND_2636 = {1{`RANDOM}};
  r_2667 = _RAND_2636[0:0];
  _RAND_2637 = {1{`RANDOM}};
  r_2668 = _RAND_2637[0:0];
  _RAND_2638 = {1{`RANDOM}};
  r_2669 = _RAND_2638[0:0];
  _RAND_2639 = {1{`RANDOM}};
  r_2670 = _RAND_2639[0:0];
  _RAND_2640 = {1{`RANDOM}};
  r_2671 = _RAND_2640[0:0];
  _RAND_2641 = {1{`RANDOM}};
  r_2672 = _RAND_2641[0:0];
  _RAND_2642 = {1{`RANDOM}};
  r_2673 = _RAND_2642[0:0];
  _RAND_2643 = {1{`RANDOM}};
  r_2674 = _RAND_2643[0:0];
  _RAND_2644 = {1{`RANDOM}};
  r_2675 = _RAND_2644[0:0];
  _RAND_2645 = {1{`RANDOM}};
  r_2676 = _RAND_2645[0:0];
  _RAND_2646 = {1{`RANDOM}};
  r_2677 = _RAND_2646[0:0];
  _RAND_2647 = {1{`RANDOM}};
  r_2678 = _RAND_2647[0:0];
  _RAND_2648 = {1{`RANDOM}};
  r_2679 = _RAND_2648[0:0];
  _RAND_2649 = {1{`RANDOM}};
  r_2680 = _RAND_2649[0:0];
  _RAND_2650 = {1{`RANDOM}};
  r_2681 = _RAND_2650[0:0];
  _RAND_2651 = {1{`RANDOM}};
  r_2682 = _RAND_2651[0:0];
  _RAND_2652 = {1{`RANDOM}};
  r_2683 = _RAND_2652[0:0];
  _RAND_2653 = {1{`RANDOM}};
  r_2684 = _RAND_2653[0:0];
  _RAND_2654 = {1{`RANDOM}};
  r_2685 = _RAND_2654[0:0];
  _RAND_2655 = {1{`RANDOM}};
  r_2686 = _RAND_2655[0:0];
  _RAND_2656 = {1{`RANDOM}};
  r_2687 = _RAND_2656[0:0];
  _RAND_2657 = {1{`RANDOM}};
  r_2688 = _RAND_2657[0:0];
  _RAND_2658 = {1{`RANDOM}};
  r_2689 = _RAND_2658[0:0];
  _RAND_2659 = {1{`RANDOM}};
  r_2690 = _RAND_2659[0:0];
  _RAND_2660 = {1{`RANDOM}};
  r_2691 = _RAND_2660[0:0];
  _RAND_2661 = {1{`RANDOM}};
  r_2692 = _RAND_2661[0:0];
  _RAND_2662 = {1{`RANDOM}};
  r_2693 = _RAND_2662[0:0];
  _RAND_2663 = {1{`RANDOM}};
  r_2694 = _RAND_2663[0:0];
  _RAND_2664 = {1{`RANDOM}};
  r_2695 = _RAND_2664[0:0];
  _RAND_2665 = {1{`RANDOM}};
  r_2696 = _RAND_2665[0:0];
  _RAND_2666 = {1{`RANDOM}};
  r_2697 = _RAND_2666[0:0];
  _RAND_2667 = {1{`RANDOM}};
  r_2698 = _RAND_2667[0:0];
  _RAND_2668 = {1{`RANDOM}};
  r_2699 = _RAND_2668[0:0];
  _RAND_2669 = {1{`RANDOM}};
  r_2700 = _RAND_2669[0:0];
  _RAND_2670 = {1{`RANDOM}};
  r_2701 = _RAND_2670[0:0];
  _RAND_2671 = {1{`RANDOM}};
  r_2702 = _RAND_2671[0:0];
  _RAND_2672 = {1{`RANDOM}};
  r_2703 = _RAND_2672[0:0];
  _RAND_2673 = {1{`RANDOM}};
  r_2704 = _RAND_2673[0:0];
  _RAND_2674 = {1{`RANDOM}};
  r_2705 = _RAND_2674[0:0];
  _RAND_2675 = {1{`RANDOM}};
  r_2706 = _RAND_2675[0:0];
  _RAND_2676 = {1{`RANDOM}};
  r_2707 = _RAND_2676[0:0];
  _RAND_2677 = {1{`RANDOM}};
  r_2708 = _RAND_2677[0:0];
  _RAND_2678 = {1{`RANDOM}};
  r_2709 = _RAND_2678[0:0];
  _RAND_2679 = {1{`RANDOM}};
  r_2710 = _RAND_2679[0:0];
  _RAND_2680 = {1{`RANDOM}};
  r_2711 = _RAND_2680[0:0];
  _RAND_2681 = {1{`RANDOM}};
  r_2712 = _RAND_2681[0:0];
  _RAND_2682 = {1{`RANDOM}};
  r_2713 = _RAND_2682[0:0];
  _RAND_2683 = {1{`RANDOM}};
  r_2714 = _RAND_2683[0:0];
  _RAND_2684 = {1{`RANDOM}};
  r_2715 = _RAND_2684[0:0];
  _RAND_2685 = {1{`RANDOM}};
  r_2716 = _RAND_2685[0:0];
  _RAND_2686 = {1{`RANDOM}};
  r_2717 = _RAND_2686[0:0];
  _RAND_2687 = {1{`RANDOM}};
  r_2718 = _RAND_2687[0:0];
  _RAND_2688 = {1{`RANDOM}};
  r_2719 = _RAND_2688[0:0];
  _RAND_2689 = {1{`RANDOM}};
  r_2720 = _RAND_2689[0:0];
  _RAND_2690 = {1{`RANDOM}};
  r_2721 = _RAND_2690[0:0];
  _RAND_2691 = {1{`RANDOM}};
  r_2722 = _RAND_2691[0:0];
  _RAND_2692 = {1{`RANDOM}};
  r_2723 = _RAND_2692[0:0];
  _RAND_2693 = {1{`RANDOM}};
  r_2724 = _RAND_2693[0:0];
  _RAND_2694 = {1{`RANDOM}};
  r_2725 = _RAND_2694[0:0];
  _RAND_2695 = {1{`RANDOM}};
  r_2726 = _RAND_2695[0:0];
  _RAND_2696 = {1{`RANDOM}};
  r_2727 = _RAND_2696[0:0];
  _RAND_2697 = {1{`RANDOM}};
  r_2728 = _RAND_2697[0:0];
  _RAND_2698 = {1{`RANDOM}};
  r_2729 = _RAND_2698[0:0];
  _RAND_2699 = {1{`RANDOM}};
  r_2730 = _RAND_2699[0:0];
  _RAND_2700 = {1{`RANDOM}};
  r_2731 = _RAND_2700[0:0];
  _RAND_2701 = {1{`RANDOM}};
  r_2732 = _RAND_2701[0:0];
  _RAND_2702 = {1{`RANDOM}};
  r_2733 = _RAND_2702[0:0];
  _RAND_2703 = {1{`RANDOM}};
  r_2734 = _RAND_2703[0:0];
  _RAND_2704 = {1{`RANDOM}};
  r_2735 = _RAND_2704[0:0];
  _RAND_2705 = {1{`RANDOM}};
  r_2736 = _RAND_2705[0:0];
  _RAND_2706 = {1{`RANDOM}};
  r_2737 = _RAND_2706[0:0];
  _RAND_2707 = {1{`RANDOM}};
  r_2738 = _RAND_2707[0:0];
  _RAND_2708 = {1{`RANDOM}};
  r_2739 = _RAND_2708[0:0];
  _RAND_2709 = {1{`RANDOM}};
  r_2740 = _RAND_2709[0:0];
  _RAND_2710 = {1{`RANDOM}};
  r_2741 = _RAND_2710[0:0];
  _RAND_2711 = {1{`RANDOM}};
  r_2742 = _RAND_2711[0:0];
  _RAND_2712 = {1{`RANDOM}};
  r_2743 = _RAND_2712[0:0];
  _RAND_2713 = {1{`RANDOM}};
  r_2744 = _RAND_2713[0:0];
  _RAND_2714 = {1{`RANDOM}};
  r_2745 = _RAND_2714[0:0];
  _RAND_2715 = {1{`RANDOM}};
  r_2746 = _RAND_2715[0:0];
  _RAND_2716 = {1{`RANDOM}};
  r_2747 = _RAND_2716[0:0];
  _RAND_2717 = {1{`RANDOM}};
  r_2748 = _RAND_2717[0:0];
  _RAND_2718 = {1{`RANDOM}};
  r_2749 = _RAND_2718[0:0];
  _RAND_2719 = {1{`RANDOM}};
  r_2750 = _RAND_2719[0:0];
  _RAND_2720 = {1{`RANDOM}};
  r_2751 = _RAND_2720[0:0];
  _RAND_2721 = {1{`RANDOM}};
  r_2752 = _RAND_2721[0:0];
  _RAND_2722 = {1{`RANDOM}};
  r_2753 = _RAND_2722[0:0];
  _RAND_2723 = {1{`RANDOM}};
  r_2754 = _RAND_2723[0:0];
  _RAND_2724 = {1{`RANDOM}};
  r_2755 = _RAND_2724[0:0];
  _RAND_2725 = {1{`RANDOM}};
  r_2756 = _RAND_2725[0:0];
  _RAND_2726 = {1{`RANDOM}};
  r_2757 = _RAND_2726[0:0];
  _RAND_2727 = {1{`RANDOM}};
  r_2758 = _RAND_2727[0:0];
  _RAND_2728 = {1{`RANDOM}};
  r_2759 = _RAND_2728[0:0];
  _RAND_2729 = {1{`RANDOM}};
  r_2760 = _RAND_2729[0:0];
  _RAND_2730 = {1{`RANDOM}};
  r_2761 = _RAND_2730[0:0];
  _RAND_2731 = {1{`RANDOM}};
  r_2762 = _RAND_2731[0:0];
  _RAND_2732 = {1{`RANDOM}};
  r_2763 = _RAND_2732[0:0];
  _RAND_2733 = {1{`RANDOM}};
  r_2764 = _RAND_2733[0:0];
  _RAND_2734 = {1{`RANDOM}};
  r_2765 = _RAND_2734[0:0];
  _RAND_2735 = {1{`RANDOM}};
  r_2766 = _RAND_2735[0:0];
  _RAND_2736 = {1{`RANDOM}};
  r_2767 = _RAND_2736[0:0];
  _RAND_2737 = {1{`RANDOM}};
  r_2768 = _RAND_2737[0:0];
  _RAND_2738 = {1{`RANDOM}};
  r_2769 = _RAND_2738[0:0];
  _RAND_2739 = {1{`RANDOM}};
  r_2770 = _RAND_2739[0:0];
  _RAND_2740 = {1{`RANDOM}};
  r_2771 = _RAND_2740[0:0];
  _RAND_2741 = {1{`RANDOM}};
  r_2772 = _RAND_2741[0:0];
  _RAND_2742 = {1{`RANDOM}};
  r_2773 = _RAND_2742[0:0];
  _RAND_2743 = {1{`RANDOM}};
  r_2774 = _RAND_2743[0:0];
  _RAND_2744 = {1{`RANDOM}};
  r_2775 = _RAND_2744[0:0];
  _RAND_2745 = {1{`RANDOM}};
  r_2776 = _RAND_2745[0:0];
  _RAND_2746 = {1{`RANDOM}};
  r_2777 = _RAND_2746[0:0];
  _RAND_2747 = {1{`RANDOM}};
  r_2778 = _RAND_2747[0:0];
  _RAND_2748 = {1{`RANDOM}};
  r_2779 = _RAND_2748[0:0];
  _RAND_2749 = {1{`RANDOM}};
  r_2780 = _RAND_2749[0:0];
  _RAND_2750 = {1{`RANDOM}};
  r_2781 = _RAND_2750[0:0];
  _RAND_2751 = {1{`RANDOM}};
  r_2782 = _RAND_2751[0:0];
  _RAND_2752 = {1{`RANDOM}};
  r_2783 = _RAND_2752[0:0];
  _RAND_2753 = {1{`RANDOM}};
  r_2784 = _RAND_2753[0:0];
  _RAND_2754 = {1{`RANDOM}};
  r_2785 = _RAND_2754[0:0];
  _RAND_2755 = {1{`RANDOM}};
  r_2786 = _RAND_2755[0:0];
  _RAND_2756 = {1{`RANDOM}};
  r_2787 = _RAND_2756[0:0];
  _RAND_2757 = {1{`RANDOM}};
  r_2788 = _RAND_2757[0:0];
  _RAND_2758 = {1{`RANDOM}};
  r_2789 = _RAND_2758[0:0];
  _RAND_2759 = {1{`RANDOM}};
  r_2790 = _RAND_2759[0:0];
  _RAND_2760 = {1{`RANDOM}};
  r_2791 = _RAND_2760[0:0];
  _RAND_2761 = {1{`RANDOM}};
  r_2792 = _RAND_2761[0:0];
  _RAND_2762 = {1{`RANDOM}};
  r_2793 = _RAND_2762[0:0];
  _RAND_2763 = {1{`RANDOM}};
  r_2794 = _RAND_2763[0:0];
  _RAND_2764 = {1{`RANDOM}};
  r_2795 = _RAND_2764[0:0];
  _RAND_2765 = {1{`RANDOM}};
  r_2796 = _RAND_2765[0:0];
  _RAND_2766 = {1{`RANDOM}};
  r_2797 = _RAND_2766[0:0];
  _RAND_2767 = {1{`RANDOM}};
  r_2798 = _RAND_2767[0:0];
  _RAND_2768 = {1{`RANDOM}};
  r_2799 = _RAND_2768[0:0];
  _RAND_2769 = {1{`RANDOM}};
  r_2800 = _RAND_2769[0:0];
  _RAND_2770 = {1{`RANDOM}};
  r_2801 = _RAND_2770[0:0];
  _RAND_2771 = {1{`RANDOM}};
  r_2802 = _RAND_2771[0:0];
  _RAND_2772 = {1{`RANDOM}};
  r_2803 = _RAND_2772[0:0];
  _RAND_2773 = {1{`RANDOM}};
  r_2804 = _RAND_2773[0:0];
  _RAND_2774 = {1{`RANDOM}};
  r_2805 = _RAND_2774[0:0];
  _RAND_2775 = {1{`RANDOM}};
  r_2806 = _RAND_2775[0:0];
  _RAND_2776 = {1{`RANDOM}};
  r_2807 = _RAND_2776[0:0];
  _RAND_2777 = {1{`RANDOM}};
  r_2808 = _RAND_2777[0:0];
  _RAND_2778 = {1{`RANDOM}};
  r_2809 = _RAND_2778[0:0];
  _RAND_2779 = {1{`RANDOM}};
  r_2810 = _RAND_2779[0:0];
  _RAND_2780 = {1{`RANDOM}};
  r_2811 = _RAND_2780[0:0];
  _RAND_2781 = {1{`RANDOM}};
  r_2812 = _RAND_2781[0:0];
  _RAND_2782 = {1{`RANDOM}};
  r_2813 = _RAND_2782[0:0];
  _RAND_2783 = {1{`RANDOM}};
  r_2814 = _RAND_2783[0:0];
  _RAND_2784 = {1{`RANDOM}};
  r_2815 = _RAND_2784[0:0];
  _RAND_2785 = {1{`RANDOM}};
  r_2816 = _RAND_2785[0:0];
  _RAND_2786 = {1{`RANDOM}};
  r_2817 = _RAND_2786[0:0];
  _RAND_2787 = {1{`RANDOM}};
  r_2818 = _RAND_2787[0:0];
  _RAND_2788 = {1{`RANDOM}};
  r_2819 = _RAND_2788[0:0];
  _RAND_2789 = {1{`RANDOM}};
  r_2820 = _RAND_2789[0:0];
  _RAND_2790 = {1{`RANDOM}};
  r_2821 = _RAND_2790[0:0];
  _RAND_2791 = {1{`RANDOM}};
  r_2822 = _RAND_2791[0:0];
  _RAND_2792 = {1{`RANDOM}};
  r_2823 = _RAND_2792[0:0];
  _RAND_2793 = {1{`RANDOM}};
  r_2824 = _RAND_2793[0:0];
  _RAND_2794 = {1{`RANDOM}};
  r_2825 = _RAND_2794[0:0];
  _RAND_2795 = {1{`RANDOM}};
  r_2826 = _RAND_2795[0:0];
  _RAND_2796 = {1{`RANDOM}};
  r_2827 = _RAND_2796[0:0];
  _RAND_2797 = {1{`RANDOM}};
  r_2828 = _RAND_2797[0:0];
  _RAND_2798 = {1{`RANDOM}};
  r_2829 = _RAND_2798[0:0];
  _RAND_2799 = {1{`RANDOM}};
  r_2830 = _RAND_2799[0:0];
  _RAND_2800 = {1{`RANDOM}};
  r_2831 = _RAND_2800[0:0];
  _RAND_2801 = {1{`RANDOM}};
  r_2832 = _RAND_2801[0:0];
  _RAND_2802 = {1{`RANDOM}};
  r_2833 = _RAND_2802[0:0];
  _RAND_2803 = {1{`RANDOM}};
  r_2834 = _RAND_2803[0:0];
  _RAND_2804 = {1{`RANDOM}};
  r_2835 = _RAND_2804[0:0];
  _RAND_2805 = {1{`RANDOM}};
  r_2836 = _RAND_2805[0:0];
  _RAND_2806 = {1{`RANDOM}};
  r_2837 = _RAND_2806[0:0];
  _RAND_2807 = {1{`RANDOM}};
  r_2838 = _RAND_2807[0:0];
  _RAND_2808 = {1{`RANDOM}};
  r_2839 = _RAND_2808[0:0];
  _RAND_2809 = {1{`RANDOM}};
  r_2840 = _RAND_2809[0:0];
  _RAND_2810 = {1{`RANDOM}};
  r_2841 = _RAND_2810[0:0];
  _RAND_2811 = {1{`RANDOM}};
  r_2842 = _RAND_2811[0:0];
  _RAND_2812 = {1{`RANDOM}};
  r_2843 = _RAND_2812[0:0];
  _RAND_2813 = {1{`RANDOM}};
  r_2844 = _RAND_2813[0:0];
  _RAND_2814 = {1{`RANDOM}};
  r_2845 = _RAND_2814[0:0];
  _RAND_2815 = {1{`RANDOM}};
  r_2846 = _RAND_2815[0:0];
  _RAND_2816 = {1{`RANDOM}};
  r_2847 = _RAND_2816[0:0];
  _RAND_2817 = {1{`RANDOM}};
  r_2848 = _RAND_2817[0:0];
  _RAND_2818 = {1{`RANDOM}};
  r_2849 = _RAND_2818[0:0];
  _RAND_2819 = {1{`RANDOM}};
  r_2850 = _RAND_2819[0:0];
  _RAND_2820 = {1{`RANDOM}};
  r_2851 = _RAND_2820[0:0];
  _RAND_2821 = {1{`RANDOM}};
  r_2852 = _RAND_2821[0:0];
  _RAND_2822 = {1{`RANDOM}};
  r_2853 = _RAND_2822[0:0];
  _RAND_2823 = {1{`RANDOM}};
  r_2854 = _RAND_2823[0:0];
  _RAND_2824 = {1{`RANDOM}};
  r_2855 = _RAND_2824[0:0];
  _RAND_2825 = {1{`RANDOM}};
  r_2856 = _RAND_2825[0:0];
  _RAND_2826 = {1{`RANDOM}};
  r_2857 = _RAND_2826[0:0];
  _RAND_2827 = {1{`RANDOM}};
  r_2858 = _RAND_2827[0:0];
  _RAND_2828 = {1{`RANDOM}};
  r_2859 = _RAND_2828[0:0];
  _RAND_2829 = {1{`RANDOM}};
  r_2860 = _RAND_2829[0:0];
  _RAND_2830 = {1{`RANDOM}};
  r_2861 = _RAND_2830[0:0];
  _RAND_2831 = {1{`RANDOM}};
  r_2862 = _RAND_2831[0:0];
  _RAND_2832 = {1{`RANDOM}};
  r_2863 = _RAND_2832[0:0];
  _RAND_2833 = {1{`RANDOM}};
  r_2864 = _RAND_2833[0:0];
  _RAND_2834 = {1{`RANDOM}};
  r_2865 = _RAND_2834[0:0];
  _RAND_2835 = {1{`RANDOM}};
  r_2866 = _RAND_2835[0:0];
  _RAND_2836 = {1{`RANDOM}};
  r_2867 = _RAND_2836[0:0];
  _RAND_2837 = {1{`RANDOM}};
  r_2868 = _RAND_2837[0:0];
  _RAND_2838 = {1{`RANDOM}};
  r_2869 = _RAND_2838[0:0];
  _RAND_2839 = {1{`RANDOM}};
  r_2870 = _RAND_2839[0:0];
  _RAND_2840 = {1{`RANDOM}};
  count = _RAND_2840[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MUL(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [63:0] io_in_bits_ctrl_data_src1,
  input  [63:0] io_in_bits_ctrl_data_src2,
  output        io_out_valid,
  output [63:0] io_out_bits_result_result_lo
);
  wire  mult_clock; // @[MUL.scala 362:24]
  wire  mult_reset; // @[MUL.scala 362:24]
  wire  mult_io_in_valid; // @[MUL.scala 362:24]
  wire [63:0] mult_io_in_bits_ctrl_data_src1; // @[MUL.scala 362:24]
  wire [63:0] mult_io_in_bits_ctrl_data_src2; // @[MUL.scala 362:24]
  wire  mult_io_out_valid; // @[MUL.scala 362:24]
  wire [63:0] mult_io_out_bits_result_result_lo; // @[MUL.scala 362:24]
  Booth_Walloc_MUL mult ( // @[MUL.scala 362:24]
    .clock(mult_clock),
    .reset(mult_reset),
    .io_in_valid(mult_io_in_valid),
    .io_in_bits_ctrl_data_src1(mult_io_in_bits_ctrl_data_src1),
    .io_in_bits_ctrl_data_src2(mult_io_in_bits_ctrl_data_src2),
    .io_out_valid(mult_io_out_valid),
    .io_out_bits_result_result_lo(mult_io_out_bits_result_result_lo)
  );
  assign io_out_valid = mult_io_out_valid; // @[MUL.scala 364:14]
  assign io_out_bits_result_result_lo = mult_io_out_bits_result_result_lo; // @[MUL.scala 364:14]
  assign mult_clock = clock;
  assign mult_reset = reset;
  assign mult_io_in_valid = io_in_valid; // @[MUL.scala 363:13]
  assign mult_io_in_bits_ctrl_data_src1 = io_in_bits_ctrl_data_src1; // @[MUL.scala 363:13]
  assign mult_io_in_bits_ctrl_data_src2 = io_in_bits_ctrl_data_src2; // @[MUL.scala 363:13]
endmodule
module DIV(
  input         clock,
  input         reset,
  input         io_in_valid,
  input         io_in_bits_ctrl_flow_div_signed,
  input  [63:0] io_in_bits_ctrl_data_src1,
  input  [63:0] io_in_bits_ctrl_data_src2,
  output        io_out_valid,
  output [63:0] io_out_bits_result_quotient,
  output [63:0] io_out_bits_result_remainder
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] dividend; // @[DIV.scala 15:25]
  reg [63:0] divisor; // @[DIV.scala 16:24]
  reg [63:0] S; // @[DIV.scala 17:18]
  reg [1:0] state; // @[DIV.scala 23:22]
  wire  _T = state == 2'h1; // @[DIV.scala 24:33]
  reg [5:0] count; // @[Counter.scala 62:40]
  wire  wrap_wrap = count == 6'h3f; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = count + 6'h1; // @[Counter.scala 78:24]
  wire  s = _T & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire [64:0] _res_div_T_1 = {1'h0,divisor}; // @[Cat.scala 31:58]
  wire [64:0] res_div = dividend[127:63] - _res_div_T_1; // @[DIV.scala 25:49]
  wire [1:0] _GEN_2 = state == 2'h0 ? 2'h1 : state; // @[DIV.scala 27:25 28:13 23:22]
  wire [63:0] _dividend_T_4 = 64'h0 - io_in_bits_ctrl_data_src1; // @[DIV.scala 43:87]
  wire [63:0] _dividend_T_5 = io_in_bits_ctrl_flow_div_signed & io_in_bits_ctrl_data_src1[63] ? _dividend_T_4 :
    io_in_bits_ctrl_data_src1; // @[DIV.scala 43:12]
  wire [127:0] _dividend_T_6 = {64'h0,_dividend_T_5}; // @[Cat.scala 31:58]
  wire [63:0] _divisor_T_3 = 64'h0 - io_in_bits_ctrl_data_src2; // @[DIV.scala 44:96]
  wire  _S_T_1 = ~res_div[64]; // @[DIV.scala 48:35]
  wire [63:0] _S_T_3 = {S[63:1],1'h1}; // @[Cat.scala 31:58]
  wire [63:0] _S_T_5 = {S[63:1],1'h0}; // @[Cat.scala 31:58]
  wire [63:0] _S_T_6 = ~res_div[64] ? _S_T_3 : _S_T_5; // @[DIV.scala 48:17]
  wire [64:0] _S_T_7 = {_S_T_6, 1'h0}; // @[DIV.scala 49:79]
  wire [64:0] _GEN_6 = count != 6'h3f ? _S_T_7 : {{1'd0}, _S_T_6}; // @[DIV.scala 47:36 48:11 51:11]
  wire [127:0] _dividend_T_14 = {res_div,dividend[62:0]}; // @[Cat.scala 31:58]
  wire [127:0] _dividend_T_15 = _S_T_1 ? _dividend_T_14 : dividend; // @[DIV.scala 54:22]
  wire [128:0] _dividend_T_16 = {_dividend_T_15, 1'h0}; // @[DIV.scala 55:110]
  wire [64:0] _GEN_7 = 2'h1 == state ? _GEN_6 : {{1'd0}, S}; // @[DIV.scala 40:16 17:18]
  wire [128:0] _GEN_8 = 2'h1 == state ? _dividend_T_16 : {{1'd0}, dividend}; // @[DIV.scala 40:16 54:16 15:25]
  wire [128:0] _GEN_9 = 2'h0 == state ? {{1'd0}, _dividend_T_6} : _GEN_8; // @[DIV.scala 40:16 42:16]
  wire [64:0] _GEN_11 = 2'h0 == state ? {{1'd0}, S} : _GEN_7; // @[DIV.scala 40:16 17:18]
  wire [63:0] negative_s = 64'h0 - S; // @[DIV.scala 63:20]
  wire [63:0] negative_r = 64'h0 - dividend[127:64]; // @[DIV.scala 64:20]
  wire [63:0] _T_13 = S[63] ? negative_s : S; // @[DIV.scala 67:18]
  wire [63:0] _T_16 = dividend[127] ? negative_r : dividend[127:64]; // @[DIV.scala 67:49]
  wire [63:0] _T_18 = S[63] ? S : negative_s; // @[DIV.scala 68:18]
  wire [63:0] _T_26 = dividend[127] ? dividend[127:64] : negative_r; // @[DIV.scala 69:49]
  wire [1:0] _s_o_T_2 = {io_in_bits_ctrl_data_src1[63],io_in_bits_ctrl_data_src2[63]}; // @[Cat.scala 31:58]
  wire  _s_o_T_3 = 2'h0 == _s_o_T_2; // @[util.scala 45:32]
  wire  _s_o_T_4 = 2'h1 == _s_o_T_2; // @[util.scala 45:32]
  wire  _s_o_T_5 = 2'h2 == _s_o_T_2; // @[util.scala 45:32]
  wire  _s_o_T_6 = 2'h3 == _s_o_T_2; // @[util.scala 45:32]
  wire [63:0] _s_o_T_7 = _s_o_T_3 ? _T_13 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _s_o_T_8 = _s_o_T_4 ? _T_18 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _s_o_T_9 = _s_o_T_5 ? _T_18 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _s_o_T_10 = _s_o_T_6 ? _T_13 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _s_o_T_11 = _s_o_T_7 | _s_o_T_8; // @[Mux.scala 27:73]
  wire [63:0] _s_o_T_12 = _s_o_T_11 | _s_o_T_9; // @[Mux.scala 27:73]
  wire [63:0] s_o = _s_o_T_12 | _s_o_T_10; // @[Mux.scala 27:73]
  wire [63:0] _r_o_T_7 = _s_o_T_3 ? _T_16 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _r_o_T_8 = _s_o_T_4 ? _T_16 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _r_o_T_9 = _s_o_T_5 ? _T_26 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _r_o_T_10 = _s_o_T_6 ? _T_26 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _r_o_T_11 = _r_o_T_7 | _r_o_T_8; // @[Mux.scala 27:73]
  wire [63:0] _r_o_T_12 = _r_o_T_11 | _r_o_T_9; // @[Mux.scala 27:73]
  wire [63:0] r_o = _r_o_T_12 | _r_o_T_10; // @[Mux.scala 27:73]
  wire [128:0] _GEN_12 = reset ? 129'h0 : _GEN_9; // @[DIV.scala 15:{25,25}]
  wire [64:0] _GEN_13 = reset ? 65'h0 : _GEN_11; // @[DIV.scala 17:{18,18}]
  assign io_out_valid = state == 2'h2; // @[DIV.scala 76:29]
  assign io_out_bits_result_quotient = io_in_bits_ctrl_flow_div_signed ? s_o : S; // @[DIV.scala 77:37]
  assign io_out_bits_result_remainder = io_in_bits_ctrl_flow_div_signed ? r_o : dividend[127:64]; // @[DIV.scala 78:38]
  always @(posedge clock) begin
    dividend <= _GEN_12[127:0]; // @[DIV.scala 15:{25,25}]
    if (reset) begin // @[DIV.scala 16:24]
      divisor <= 64'h0; // @[DIV.scala 16:24]
    end else if (2'h0 == state) begin // @[DIV.scala 40:16]
      if (io_in_bits_ctrl_flow_div_signed & io_in_bits_ctrl_data_src2[63]) begin // @[DIV.scala 44:21]
        divisor <= _divisor_T_3;
      end else begin
        divisor <= io_in_bits_ctrl_data_src2;
      end
    end
    S <= _GEN_13[63:0]; // @[DIV.scala 17:{18,18}]
    if (reset) begin // @[DIV.scala 23:22]
      state <= 2'h0; // @[DIV.scala 23:22]
    end else if (io_in_valid) begin // @[DIV.scala 26:51]
      if (state == 2'h2) begin // @[DIV.scala 33:24]
        state <= 2'h0; // @[DIV.scala 34:13]
      end else if (_T & s) begin // @[DIV.scala 30:40]
        state <= 2'h2; // @[DIV.scala 31:15]
      end else begin
        state <= _GEN_2;
      end
    end else begin
      state <= 2'h0; // @[DIV.scala 37:11]
    end
    if (reset) begin // @[Counter.scala 62:40]
      count <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T) begin // @[Counter.scala 120:16]
      count <= _wrap_value_T_1; // @[Counter.scala 78:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  dividend = _RAND_0[127:0];
  _RAND_1 = {2{`RANDOM}};
  divisor = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  S = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  count = _RAND_4[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EXE(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [2:0]  io_in_bits_ctrl_signal_src1Type,
  input  [2:0]  io_in_bits_ctrl_signal_src2Type,
  input  [2:0]  io_in_bits_ctrl_signal_fuType,
  input         io_in_bits_ctrl_signal_inst_valid,
  input  [4:0]  io_in_bits_ctrl_signal_rfSrc1,
  input  [4:0]  io_in_bits_ctrl_signal_rfSrc2,
  input         io_in_bits_ctrl_signal_rfWen,
  input  [6:0]  io_in_bits_ctrl_signal_aluoptype,
  input  [4:0]  io_in_bits_ctrl_signal_rfDest,
  input  [63:0] io_in_bits_ctrl_data_src1,
  input  [63:0] io_in_bits_ctrl_data_src2,
  input  [63:0] io_in_bits_ctrl_data_Imm,
  input  [63:0] io_in_bits_ctrl_flow_PC,
  input  [31:0] io_in_bits_ctrl_flow_inst,
  input  [63:0] io_src1,
  input  [63:0] io_src2,
  output        io_branchIO_is_branch,
  output        io_branchIO_is_jump,
  output [63:0] io_branchIO_dnpc,
  input         io_out_ready,
  output        io_out_valid,
  output [2:0]  io_out_bits_ctrl_signal_fuType,
  output        io_out_bits_ctrl_signal_inst_valid,
  output        io_out_bits_ctrl_signal_rfWen,
  output [6:0]  io_out_bits_ctrl_signal_aluoptype,
  output [63:0] io_out_bits_ctrl_flow_PC,
  output [31:0] io_out_bits_ctrl_flow_inst,
  output [63:0] io_out_bits_ctrl_flow_Dnpc,
  output [4:0]  io_out_bits_ctrl_rf_rfDest,
  output        io_out_bits_ctrl_rf_rfWen,
  output [63:0] io_out_bits_ctrl_rf_rfData,
  output [63:0] io_out_bits_ctrl_data_src1,
  output [63:0] io_out_bits_ctrl_data_src2,
  output [63:0] io_out_bits_ctrl_data_Imm,
  output        io_is_break,
  output        io_is_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] CSRDIFF_mepc; // @[EXE.scala 115:21]
  wire [63:0] CSRDIFF_mcause; // @[EXE.scala 115:21]
  wire [63:0] CSRDIFF_mstatus; // @[EXE.scala 115:21]
  wire [63:0] CSRDIFF_mtvec; // @[EXE.scala 115:21]
  wire  mul_clock; // @[EXE.scala 118:19]
  wire  mul_reset; // @[EXE.scala 118:19]
  wire  mul_io_in_valid; // @[EXE.scala 118:19]
  wire [63:0] mul_io_in_bits_ctrl_data_src1; // @[EXE.scala 118:19]
  wire [63:0] mul_io_in_bits_ctrl_data_src2; // @[EXE.scala 118:19]
  wire  mul_io_out_valid; // @[EXE.scala 118:19]
  wire [63:0] mul_io_out_bits_result_result_lo; // @[EXE.scala 118:19]
  wire  div_clock; // @[EXE.scala 119:19]
  wire  div_reset; // @[EXE.scala 119:19]
  wire  div_io_in_valid; // @[EXE.scala 119:19]
  wire  div_io_in_bits_ctrl_flow_div_signed; // @[EXE.scala 119:19]
  wire [63:0] div_io_in_bits_ctrl_data_src1; // @[EXE.scala 119:19]
  wire [63:0] div_io_in_bits_ctrl_data_src2; // @[EXE.scala 119:19]
  wire  div_io_out_valid; // @[EXE.scala 119:19]
  wire [63:0] div_io_out_bits_result_quotient; // @[EXE.scala 119:19]
  wire [63:0] div_io_out_bits_result_remainder; // @[EXE.scala 119:19]
  wire  _is_mul_T = 7'h78 == io_in_bits_ctrl_signal_aluoptype; // @[EXE.scala 104:32]
  wire  _is_mul_T_1 = 7'h7 == io_in_bits_ctrl_signal_aluoptype; // @[EXE.scala 104:86]
  wire  is_mul = (7'h78 == io_in_bits_ctrl_signal_aluoptype | 7'h7 == io_in_bits_ctrl_signal_aluoptype) &
    io_in_bits_ctrl_signal_inst_valid & io_in_valid; // @[EXE.scala 104:161]
  wire  _is_div_T = io_in_bits_ctrl_signal_aluoptype == 7'h43; // @[EXE.scala 105:50]
  wire  _is_div_T_2 = io_in_bits_ctrl_signal_aluoptype == 7'h43 | io_in_bits_ctrl_signal_aluoptype == 7'h13; // @[EXE.scala 105:68]
  wire  _is_div_T_3 = io_in_bits_ctrl_signal_aluoptype == 7'h79; // @[EXE.scala 106:41]
  wire  _is_div_T_5 = io_in_bits_ctrl_signal_aluoptype == 7'h10; // @[EXE.scala 106:96]
  wire  _is_div_T_6 = _is_div_T_2 | io_in_bits_ctrl_signal_aluoptype == 7'h79 | io_in_bits_ctrl_signal_aluoptype == 7'h10
    ; // @[EXE.scala 106:60]
  wire  _is_div_T_7 = io_in_bits_ctrl_signal_aluoptype == 7'h12; // @[EXE.scala 107:41]
  wire  _is_div_T_10 = _is_div_T_6 | io_in_bits_ctrl_signal_aluoptype == 7'h12 | io_in_bits_ctrl_signal_aluoptype == 7'hf
    ; // @[EXE.scala 107:59]
  wire  _is_div_T_11 = io_in_bits_ctrl_signal_aluoptype == 7'h7a; // @[EXE.scala 108:41]
  wire  _is_div_T_13 = io_in_bits_ctrl_signal_aluoptype == 7'hd; // @[EXE.scala 108:96]
  wire  is_div = (_is_div_T_10 | io_in_bits_ctrl_signal_aluoptype == 7'h7a | io_in_bits_ctrl_signal_aluoptype == 7'hd)
     & io_in_bits_ctrl_signal_inst_valid & io_in_valid; // @[EXE.scala 108:154]
  wire  _is_divw_T_2 = _is_div_T_3 | _is_div_T_5; // @[EXE.scala 109:70]
  wire  is_divw = _is_divw_T_2 | _is_div_T_11 | _is_div_T_13; // @[EXE.scala 110:60]
  wire  _is_div_sign_T_2 = _is_div_T | _is_div_T_3; // @[EXE.scala 111:73]
  wire  is_div_sign = _is_div_sign_T_2 | _is_div_T_7 | _is_div_T_11; // @[EXE.scala 112:59]
  reg [63:0] mepc; // @[CSR.scala 18:17]
  reg [63:0] mcause; // @[CSR.scala 19:23]
  reg [63:0] mstatus; // @[CSR.scala 20:24]
  reg [63:0] mtvec; // @[CSR.scala 21:22]
  reg [63:0] mie; // @[CSR.scala 22:20]
  reg [63:0] mip; // @[CSR.scala 23:20]
  wire [63:0] _GEN_1 = 3'h2 == io_in_bits_ctrl_signal_src1Type ? io_in_bits_ctrl_flow_PC : 64'h0; // @[EXE.scala 124:43 129:12]
  wire [63:0] src1 = 3'h0 == io_in_bits_ctrl_signal_src1Type ? io_src1 : _GEN_1; // @[EXE.scala 124:43 126:12]
  wire [63:0] _GEN_3 = 3'h1 == io_in_bits_ctrl_signal_src2Type ? io_in_bits_ctrl_data_Imm : 64'h0; // @[EXE.scala 135:43 141:12]
  wire [63:0] src2 = 3'h0 == io_in_bits_ctrl_signal_src2Type ? io_src2 : _GEN_3; // @[EXE.scala 135:43 138:12]
  wire [63:0] _dnpc_T_1 = io_in_bits_ctrl_flow_PC + 64'h4; // @[EXE.scala 147:49]
  wire [63:0] _alu_result_T_1 = src1 + src2; // @[EXE.scala 158:26]
  wire  alu_result_sign = _alu_result_T_1[31]; // @[util.scala 11:19]
  wire [31:0] _alu_result_T_6 = alu_result_sign ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_result_T_7 = {_alu_result_T_6,_alu_result_T_1[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _alu_result_T_8 = src1 | src2; // @[EXE.scala 167:26]
  wire [63:0] _alu_result_T_10 = src1 - src2; // @[EXE.scala 170:26]
  wire [63:0] _alu_result_T_11 = src1 & src2; // @[EXE.scala 173:26]
  wire [63:0] _alu_result_T_12 = src1 ^ src2; // @[EXE.scala 176:26]
  wire  alu_result_sign_2 = mul_io_out_bits_result_result_lo[31]; // @[util.scala 11:19]
  wire [31:0] _alu_result_T_21 = alu_result_sign_2 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_result_T_22 = {_alu_result_T_21,mul_io_out_bits_result_result_lo[31:0]}; // @[Cat.scala 31:58]
  wire  alu_result_sign_3 = div_io_out_bits_result_quotient[31]; // @[util.scala 11:19]
  wire [31:0] _alu_result_T_25 = alu_result_sign_3 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_result_T_26 = {_alu_result_T_25,div_io_out_bits_result_quotient[31:0]}; // @[Cat.scala 31:58]
  wire  alu_result_sign_4 = div_io_out_bits_result_remainder[31]; // @[util.scala 11:19]
  wire [31:0] _alu_result_T_29 = alu_result_sign_4 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_result_T_30 = {_alu_result_T_29,div_io_out_bits_result_remainder[31:0]}; // @[Cat.scala 31:58]
  wire  alu_result_sign_6 = _alu_result_T_10[31]; // @[util.scala 11:19]
  wire [31:0] _alu_result_T_39 = alu_result_sign_6 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _alu_result_T_40 = {_alu_result_T_39,_alu_result_T_10[31:0]}; // @[Cat.scala 31:58]
  wire  _alu_result_T_46 = io_in_bits_ctrl_data_Imm[11:0] == 12'h300; // @[CSR.scala 26:11]
  wire  _alu_result_T_47 = io_in_bits_ctrl_data_Imm[11:0] == 12'h305; // @[CSR.scala 27:11]
  wire  _alu_result_T_48 = io_in_bits_ctrl_data_Imm[11:0] == 12'h341; // @[CSR.scala 28:11]
  wire  _alu_result_T_49 = io_in_bits_ctrl_data_Imm[11:0] == 12'h342; // @[CSR.scala 29:11]
  wire  _alu_result_T_50 = io_in_bits_ctrl_data_Imm[11:0] == 12'h304; // @[CSR.scala 30:11]
  wire  _alu_result_T_51 = io_in_bits_ctrl_data_Imm[11:0] == 12'h344; // @[CSR.scala 31:11]
  wire [63:0] _alu_result_T_52 = _alu_result_T_51 ? mip : 64'h0; // @[Mux.scala 101:16]
  wire [63:0] _alu_result_T_53 = _alu_result_T_50 ? mie : _alu_result_T_52; // @[Mux.scala 101:16]
  wire [63:0] _alu_result_T_54 = _alu_result_T_49 ? mcause : _alu_result_T_53; // @[Mux.scala 101:16]
  wire [63:0] _alu_result_T_55 = _alu_result_T_48 ? mepc : _alu_result_T_54; // @[Mux.scala 101:16]
  wire [63:0] _alu_result_T_56 = _alu_result_T_47 ? mtvec : _alu_result_T_55; // @[Mux.scala 101:16]
  wire [63:0] _alu_result_T_57 = _alu_result_T_46 ? mstatus : _alu_result_T_56; // @[Mux.scala 101:16]
  wire [63:0] _T_39 = _alu_result_T_57 | src1; // @[EXE.scala 216:50]
  wire [63:0] _GEN_5 = _alu_result_T_51 ? _T_39 : mip; // @[CSR.scala 50:41 51:13 23:20]
  wire [63:0] _GEN_6 = _alu_result_T_50 ? _T_39 : mie; // @[CSR.scala 47:41 48:13 22:20]
  wire [63:0] _GEN_7 = _alu_result_T_50 ? mip : _GEN_5; // @[CSR.scala 23:20 47:41]
  wire [63:0] _GEN_8 = _alu_result_T_49 ? _T_39 : mcause; // @[CSR.scala 44:44 45:16 19:23]
  wire [63:0] _GEN_9 = _alu_result_T_49 ? mie : _GEN_6; // @[CSR.scala 22:20 44:44]
  wire [63:0] _GEN_10 = _alu_result_T_49 ? mip : _GEN_7; // @[CSR.scala 23:20 44:44]
  wire [63:0] _GEN_11 = _alu_result_T_48 ? _T_39 : mepc; // @[CSR.scala 41:42 42:14 18:17]
  wire [63:0] _GEN_12 = _alu_result_T_48 ? mcause : _GEN_8; // @[CSR.scala 19:23 41:42]
  wire [63:0] _GEN_13 = _alu_result_T_48 ? mie : _GEN_9; // @[CSR.scala 22:20 41:42]
  wire [63:0] _GEN_14 = _alu_result_T_48 ? mip : _GEN_10; // @[CSR.scala 23:20 41:42]
  wire [63:0] _GEN_15 = _alu_result_T_47 ? _T_39 : mtvec; // @[CSR.scala 38:43 39:15 21:22]
  wire [63:0] _GEN_16 = _alu_result_T_47 ? mepc : _GEN_11; // @[CSR.scala 18:17 38:43]
  wire [63:0] _GEN_17 = _alu_result_T_47 ? mcause : _GEN_12; // @[CSR.scala 19:23 38:43]
  wire [63:0] _GEN_18 = _alu_result_T_47 ? mie : _GEN_13; // @[CSR.scala 22:20 38:43]
  wire [63:0] _GEN_19 = _alu_result_T_47 ? mip : _GEN_14; // @[CSR.scala 23:20 38:43]
  wire [63:0] _GEN_20 = _alu_result_T_46 ? _T_39 : mstatus; // @[CSR.scala 35:38 36:15 20:24]
  wire [63:0] _GEN_21 = _alu_result_T_46 ? mtvec : _GEN_15; // @[CSR.scala 21:22 35:38]
  wire [63:0] _GEN_22 = _alu_result_T_46 ? mepc : _GEN_16; // @[CSR.scala 18:17 35:38]
  wire [63:0] _GEN_23 = _alu_result_T_46 ? mcause : _GEN_17; // @[CSR.scala 19:23 35:38]
  wire [63:0] _GEN_24 = _alu_result_T_46 ? mie : _GEN_18; // @[CSR.scala 22:20 35:38]
  wire [63:0] _GEN_25 = _alu_result_T_46 ? mip : _GEN_19; // @[CSR.scala 23:20 35:38]
  wire [63:0] _GEN_26 = _alu_result_T_51 ? src1 : mip; // @[CSR.scala 50:41 51:13 23:20]
  wire [63:0] _GEN_27 = _alu_result_T_50 ? src1 : mie; // @[CSR.scala 47:41 48:13 22:20]
  wire [63:0] _GEN_28 = _alu_result_T_50 ? mip : _GEN_26; // @[CSR.scala 23:20 47:41]
  wire [63:0] _GEN_29 = _alu_result_T_49 ? src1 : mcause; // @[CSR.scala 44:44 45:16 19:23]
  wire [63:0] _GEN_30 = _alu_result_T_49 ? mie : _GEN_27; // @[CSR.scala 22:20 44:44]
  wire [63:0] _GEN_31 = _alu_result_T_49 ? mip : _GEN_28; // @[CSR.scala 23:20 44:44]
  wire [63:0] _GEN_32 = _alu_result_T_48 ? src1 : mepc; // @[CSR.scala 41:42 42:14 18:17]
  wire [63:0] _GEN_33 = _alu_result_T_48 ? mcause : _GEN_29; // @[CSR.scala 19:23 41:42]
  wire [63:0] _GEN_34 = _alu_result_T_48 ? mie : _GEN_30; // @[CSR.scala 22:20 41:42]
  wire [63:0] _GEN_35 = _alu_result_T_48 ? mip : _GEN_31; // @[CSR.scala 23:20 41:42]
  wire [63:0] _GEN_36 = _alu_result_T_47 ? src1 : mtvec; // @[CSR.scala 38:43 39:15 21:22]
  wire [63:0] _GEN_37 = _alu_result_T_47 ? mepc : _GEN_32; // @[CSR.scala 18:17 38:43]
  wire [63:0] _GEN_38 = _alu_result_T_47 ? mcause : _GEN_33; // @[CSR.scala 19:23 38:43]
  wire [63:0] _GEN_39 = _alu_result_T_47 ? mie : _GEN_34; // @[CSR.scala 22:20 38:43]
  wire [63:0] _GEN_40 = _alu_result_T_47 ? mip : _GEN_35; // @[CSR.scala 23:20 38:43]
  wire [63:0] _GEN_41 = _alu_result_T_46 ? src1 : mstatus; // @[CSR.scala 35:38 36:15 20:24]
  wire [63:0] _GEN_42 = _alu_result_T_46 ? mtvec : _GEN_36; // @[CSR.scala 21:22 35:38]
  wire [63:0] _GEN_43 = _alu_result_T_46 ? mepc : _GEN_37; // @[CSR.scala 18:17 35:38]
  wire [63:0] _GEN_44 = _alu_result_T_46 ? mcause : _GEN_38; // @[CSR.scala 19:23 35:38]
  wire [63:0] _GEN_45 = _alu_result_T_46 ? mie : _GEN_39; // @[CSR.scala 22:20 35:38]
  wire [63:0] _GEN_46 = _alu_result_T_46 ? mip : _GEN_40; // @[CSR.scala 23:20 35:38]
  wire [63:0] _GEN_47 = 7'h16 == io_in_bits_ctrl_signal_aluoptype ? _alu_result_T_57 : 64'h0; // @[EXE.scala 156:44 219:18]
  wire [63:0] _GEN_48 = 7'h16 == io_in_bits_ctrl_signal_aluoptype ? _GEN_41 : mstatus; // @[EXE.scala 156:44 CSR.scala 20:24]
  wire [63:0] _GEN_49 = 7'h16 == io_in_bits_ctrl_signal_aluoptype ? _GEN_42 : mtvec; // @[EXE.scala 156:44 CSR.scala 21:22]
  wire [63:0] _GEN_50 = 7'h16 == io_in_bits_ctrl_signal_aluoptype ? _GEN_43 : mepc; // @[EXE.scala 156:44 CSR.scala 18:17]
  wire [63:0] _GEN_51 = 7'h16 == io_in_bits_ctrl_signal_aluoptype ? _GEN_44 : mcause; // @[EXE.scala 156:44 CSR.scala 19:23]
  wire [63:0] _GEN_52 = 7'h16 == io_in_bits_ctrl_signal_aluoptype ? _GEN_45 : mie; // @[EXE.scala 156:44 CSR.scala 22:20]
  wire [63:0] _GEN_53 = 7'h16 == io_in_bits_ctrl_signal_aluoptype ? _GEN_46 : mip; // @[EXE.scala 156:44 CSR.scala 23:20]
  wire [63:0] _GEN_54 = 7'h15 == io_in_bits_ctrl_signal_aluoptype ? _alu_result_T_57 : _GEN_47; // @[EXE.scala 156:44 215:18]
  wire [63:0] _GEN_55 = 7'h15 == io_in_bits_ctrl_signal_aluoptype ? _GEN_20 : _GEN_48; // @[EXE.scala 156:44]
  wire [63:0] _GEN_56 = 7'h15 == io_in_bits_ctrl_signal_aluoptype ? _GEN_21 : _GEN_49; // @[EXE.scala 156:44]
  wire [63:0] _GEN_57 = 7'h15 == io_in_bits_ctrl_signal_aluoptype ? _GEN_22 : _GEN_50; // @[EXE.scala 156:44]
  wire [63:0] _GEN_58 = 7'h15 == io_in_bits_ctrl_signal_aluoptype ? _GEN_23 : _GEN_51; // @[EXE.scala 156:44]
  wire [63:0] _GEN_59 = 7'h15 == io_in_bits_ctrl_signal_aluoptype ? _GEN_24 : _GEN_52; // @[EXE.scala 156:44]
  wire [63:0] _GEN_60 = 7'h15 == io_in_bits_ctrl_signal_aluoptype ? _GEN_25 : _GEN_53; // @[EXE.scala 156:44]
  wire [63:0] _GEN_61 = 7'h43 == io_in_bits_ctrl_signal_aluoptype ? div_io_out_bits_result_quotient : _GEN_54; // @[EXE.scala 156:44 212:18]
  wire [63:0] _GEN_62 = 7'h43 == io_in_bits_ctrl_signal_aluoptype ? mstatus : _GEN_55; // @[EXE.scala 156:44 CSR.scala 20:24]
  wire [63:0] _GEN_63 = 7'h43 == io_in_bits_ctrl_signal_aluoptype ? mtvec : _GEN_56; // @[EXE.scala 156:44 CSR.scala 21:22]
  wire [63:0] _GEN_64 = 7'h43 == io_in_bits_ctrl_signal_aluoptype ? mepc : _GEN_57; // @[EXE.scala 156:44 CSR.scala 18:17]
  wire [63:0] _GEN_65 = 7'h43 == io_in_bits_ctrl_signal_aluoptype ? mcause : _GEN_58; // @[EXE.scala 156:44 CSR.scala 19:23]
  wire [63:0] _GEN_66 = 7'h43 == io_in_bits_ctrl_signal_aluoptype ? mie : _GEN_59; // @[EXE.scala 156:44 CSR.scala 22:20]
  wire [63:0] _GEN_67 = 7'h43 == io_in_bits_ctrl_signal_aluoptype ? mip : _GEN_60; // @[EXE.scala 156:44 CSR.scala 23:20]
  wire [63:0] _GEN_68 = 7'h13 == io_in_bits_ctrl_signal_aluoptype ? div_io_out_bits_result_quotient : _GEN_61; // @[EXE.scala 156:44 209:18]
  wire [63:0] _GEN_69 = 7'h13 == io_in_bits_ctrl_signal_aluoptype ? mstatus : _GEN_62; // @[EXE.scala 156:44 CSR.scala 20:24]
  wire [63:0] _GEN_70 = 7'h13 == io_in_bits_ctrl_signal_aluoptype ? mtvec : _GEN_63; // @[EXE.scala 156:44 CSR.scala 21:22]
  wire [63:0] _GEN_71 = 7'h13 == io_in_bits_ctrl_signal_aluoptype ? mepc : _GEN_64; // @[EXE.scala 156:44 CSR.scala 18:17]
  wire [63:0] _GEN_72 = 7'h13 == io_in_bits_ctrl_signal_aluoptype ? mcause : _GEN_65; // @[EXE.scala 156:44 CSR.scala 19:23]
  wire [63:0] _GEN_73 = 7'h13 == io_in_bits_ctrl_signal_aluoptype ? mie : _GEN_66; // @[EXE.scala 156:44 CSR.scala 22:20]
  wire [63:0] _GEN_74 = 7'h13 == io_in_bits_ctrl_signal_aluoptype ? mip : _GEN_67; // @[EXE.scala 156:44 CSR.scala 23:20]
  wire [63:0] _GEN_75 = 7'h10 == io_in_bits_ctrl_signal_aluoptype ? _alu_result_T_26 : _GEN_68; // @[EXE.scala 156:44 206:18]
  wire [63:0] _GEN_76 = 7'h10 == io_in_bits_ctrl_signal_aluoptype ? mstatus : _GEN_69; // @[EXE.scala 156:44 CSR.scala 20:24]
  wire [63:0] _GEN_77 = 7'h10 == io_in_bits_ctrl_signal_aluoptype ? mtvec : _GEN_70; // @[EXE.scala 156:44 CSR.scala 21:22]
  wire [63:0] _GEN_78 = 7'h10 == io_in_bits_ctrl_signal_aluoptype ? mepc : _GEN_71; // @[EXE.scala 156:44 CSR.scala 18:17]
  wire [63:0] _GEN_79 = 7'h10 == io_in_bits_ctrl_signal_aluoptype ? mcause : _GEN_72; // @[EXE.scala 156:44 CSR.scala 19:23]
  wire [63:0] _GEN_80 = 7'h10 == io_in_bits_ctrl_signal_aluoptype ? mie : _GEN_73; // @[EXE.scala 156:44 CSR.scala 22:20]
  wire [63:0] _GEN_81 = 7'h10 == io_in_bits_ctrl_signal_aluoptype ? mip : _GEN_74; // @[EXE.scala 156:44 CSR.scala 23:20]
  wire [63:0] _GEN_82 = 7'h12 == io_in_bits_ctrl_signal_aluoptype ? div_io_out_bits_result_remainder : _GEN_75; // @[EXE.scala 156:44 203:18]
  wire [63:0] _GEN_83 = 7'h12 == io_in_bits_ctrl_signal_aluoptype ? mstatus : _GEN_76; // @[EXE.scala 156:44 CSR.scala 20:24]
  wire [63:0] _GEN_84 = 7'h12 == io_in_bits_ctrl_signal_aluoptype ? mtvec : _GEN_77; // @[EXE.scala 156:44 CSR.scala 21:22]
  wire [63:0] _GEN_85 = 7'h12 == io_in_bits_ctrl_signal_aluoptype ? mepc : _GEN_78; // @[EXE.scala 156:44 CSR.scala 18:17]
  wire [63:0] _GEN_86 = 7'h12 == io_in_bits_ctrl_signal_aluoptype ? mcause : _GEN_79; // @[EXE.scala 156:44 CSR.scala 19:23]
  wire [63:0] _GEN_87 = 7'h12 == io_in_bits_ctrl_signal_aluoptype ? mie : _GEN_80; // @[EXE.scala 156:44 CSR.scala 22:20]
  wire [63:0] _GEN_88 = 7'h12 == io_in_bits_ctrl_signal_aluoptype ? mip : _GEN_81; // @[EXE.scala 156:44 CSR.scala 23:20]
  wire [63:0] _GEN_89 = 7'hf == io_in_bits_ctrl_signal_aluoptype ? div_io_out_bits_result_remainder : _GEN_82; // @[EXE.scala 156:44 200:18]
  wire [63:0] _GEN_90 = 7'hf == io_in_bits_ctrl_signal_aluoptype ? mstatus : _GEN_83; // @[EXE.scala 156:44 CSR.scala 20:24]
  wire [63:0] _GEN_91 = 7'hf == io_in_bits_ctrl_signal_aluoptype ? mtvec : _GEN_84; // @[EXE.scala 156:44 CSR.scala 21:22]
  wire [63:0] _GEN_92 = 7'hf == io_in_bits_ctrl_signal_aluoptype ? mepc : _GEN_85; // @[EXE.scala 156:44 CSR.scala 18:17]
  wire [63:0] _GEN_93 = 7'hf == io_in_bits_ctrl_signal_aluoptype ? mcause : _GEN_86; // @[EXE.scala 156:44 CSR.scala 19:23]
  wire [63:0] _GEN_94 = 7'hf == io_in_bits_ctrl_signal_aluoptype ? mie : _GEN_87; // @[EXE.scala 156:44 CSR.scala 22:20]
  wire [63:0] _GEN_95 = 7'hf == io_in_bits_ctrl_signal_aluoptype ? mip : _GEN_88; // @[EXE.scala 156:44 CSR.scala 23:20]
  wire [63:0] _GEN_96 = _is_mul_T_1 ? mul_io_out_bits_result_result_lo : _GEN_89; // @[EXE.scala 156:44 197:18]
  wire [63:0] _GEN_97 = _is_mul_T_1 ? mstatus : _GEN_90; // @[EXE.scala 156:44 CSR.scala 20:24]
  wire [63:0] _GEN_98 = _is_mul_T_1 ? mtvec : _GEN_91; // @[EXE.scala 156:44 CSR.scala 21:22]
  wire [63:0] _GEN_99 = _is_mul_T_1 ? mepc : _GEN_92; // @[EXE.scala 156:44 CSR.scala 18:17]
  wire [63:0] _GEN_100 = _is_mul_T_1 ? mcause : _GEN_93; // @[EXE.scala 156:44 CSR.scala 19:23]
  wire [63:0] _GEN_101 = _is_mul_T_1 ? mie : _GEN_94; // @[EXE.scala 156:44 CSR.scala 22:20]
  wire [63:0] _GEN_102 = _is_mul_T_1 ? mip : _GEN_95; // @[EXE.scala 156:44 CSR.scala 23:20]
  wire [63:0] _GEN_103 = 7'h1 == io_in_bits_ctrl_signal_aluoptype ? _alu_result_T_40 : _GEN_96; // @[EXE.scala 156:44 194:18]
  wire [63:0] _GEN_104 = 7'h1 == io_in_bits_ctrl_signal_aluoptype ? mstatus : _GEN_97; // @[EXE.scala 156:44 CSR.scala 20:24]
  wire [63:0] _GEN_105 = 7'h1 == io_in_bits_ctrl_signal_aluoptype ? mtvec : _GEN_98; // @[EXE.scala 156:44 CSR.scala 21:22]
  wire [63:0] _GEN_106 = 7'h1 == io_in_bits_ctrl_signal_aluoptype ? mepc : _GEN_99; // @[EXE.scala 156:44 CSR.scala 18:17]
  wire [63:0] _GEN_107 = 7'h1 == io_in_bits_ctrl_signal_aluoptype ? mcause : _GEN_100; // @[EXE.scala 156:44 CSR.scala 19:23]
  wire [63:0] _GEN_108 = 7'h1 == io_in_bits_ctrl_signal_aluoptype ? mie : _GEN_101; // @[EXE.scala 156:44 CSR.scala 22:20]
  wire [63:0] _GEN_109 = 7'h1 == io_in_bits_ctrl_signal_aluoptype ? mip : _GEN_102; // @[EXE.scala 156:44 CSR.scala 23:20]
  wire [63:0] _GEN_110 = 7'hd == io_in_bits_ctrl_signal_aluoptype ? _alu_result_T_30 : _GEN_103; // @[EXE.scala 156:44 191:18]
  wire [63:0] _GEN_111 = 7'hd == io_in_bits_ctrl_signal_aluoptype ? mstatus : _GEN_104; // @[EXE.scala 156:44 CSR.scala 20:24]
  wire [63:0] _GEN_112 = 7'hd == io_in_bits_ctrl_signal_aluoptype ? mtvec : _GEN_105; // @[EXE.scala 156:44 CSR.scala 21:22]
  wire [63:0] _GEN_113 = 7'hd == io_in_bits_ctrl_signal_aluoptype ? mepc : _GEN_106; // @[EXE.scala 156:44 CSR.scala 18:17]
  wire [63:0] _GEN_114 = 7'hd == io_in_bits_ctrl_signal_aluoptype ? mcause : _GEN_107; // @[EXE.scala 156:44 CSR.scala 19:23]
  wire [63:0] _GEN_115 = 7'hd == io_in_bits_ctrl_signal_aluoptype ? mie : _GEN_108; // @[EXE.scala 156:44 CSR.scala 22:20]
  wire [63:0] _GEN_116 = 7'hd == io_in_bits_ctrl_signal_aluoptype ? mip : _GEN_109; // @[EXE.scala 156:44 CSR.scala 23:20]
  wire [63:0] _GEN_117 = 7'h7a == io_in_bits_ctrl_signal_aluoptype ? _alu_result_T_30 : _GEN_110; // @[EXE.scala 156:44 188:18]
  wire [63:0] _GEN_118 = 7'h7a == io_in_bits_ctrl_signal_aluoptype ? mstatus : _GEN_111; // @[EXE.scala 156:44 CSR.scala 20:24]
  wire [63:0] _GEN_119 = 7'h7a == io_in_bits_ctrl_signal_aluoptype ? mtvec : _GEN_112; // @[EXE.scala 156:44 CSR.scala 21:22]
  wire [63:0] _GEN_120 = 7'h7a == io_in_bits_ctrl_signal_aluoptype ? mepc : _GEN_113; // @[EXE.scala 156:44 CSR.scala 18:17]
  wire [63:0] _GEN_121 = 7'h7a == io_in_bits_ctrl_signal_aluoptype ? mcause : _GEN_114; // @[EXE.scala 156:44 CSR.scala 19:23]
  wire [63:0] _GEN_122 = 7'h7a == io_in_bits_ctrl_signal_aluoptype ? mie : _GEN_115; // @[EXE.scala 156:44 CSR.scala 22:20]
  wire [63:0] _GEN_123 = 7'h7a == io_in_bits_ctrl_signal_aluoptype ? mip : _GEN_116; // @[EXE.scala 156:44 CSR.scala 23:20]
  wire [63:0] _GEN_124 = 7'h79 == io_in_bits_ctrl_signal_aluoptype ? _alu_result_T_26 : _GEN_117; // @[EXE.scala 156:44 185:18]
  wire [63:0] _GEN_125 = 7'h79 == io_in_bits_ctrl_signal_aluoptype ? mstatus : _GEN_118; // @[EXE.scala 156:44 CSR.scala 20:24]
  wire [63:0] _GEN_126 = 7'h79 == io_in_bits_ctrl_signal_aluoptype ? mtvec : _GEN_119; // @[EXE.scala 156:44 CSR.scala 21:22]
  wire [63:0] _GEN_127 = 7'h79 == io_in_bits_ctrl_signal_aluoptype ? mepc : _GEN_120; // @[EXE.scala 156:44 CSR.scala 18:17]
  wire [63:0] _GEN_128 = 7'h79 == io_in_bits_ctrl_signal_aluoptype ? mcause : _GEN_121; // @[EXE.scala 156:44 CSR.scala 19:23]
  wire [63:0] _GEN_129 = 7'h79 == io_in_bits_ctrl_signal_aluoptype ? mie : _GEN_122; // @[EXE.scala 156:44 CSR.scala 22:20]
  wire [63:0] _GEN_130 = 7'h79 == io_in_bits_ctrl_signal_aluoptype ? mip : _GEN_123; // @[EXE.scala 156:44 CSR.scala 23:20]
  wire [63:0] _GEN_131 = _is_mul_T ? _alu_result_T_22 : _GEN_124; // @[EXE.scala 156:44 182:18]
  wire [63:0] _GEN_132 = _is_mul_T ? mstatus : _GEN_125; // @[EXE.scala 156:44 CSR.scala 20:24]
  wire [63:0] _GEN_133 = _is_mul_T ? mtvec : _GEN_126; // @[EXE.scala 156:44 CSR.scala 21:22]
  wire [63:0] _GEN_134 = _is_mul_T ? mepc : _GEN_127; // @[EXE.scala 156:44 CSR.scala 18:17]
  wire [63:0] _GEN_135 = _is_mul_T ? mcause : _GEN_128; // @[EXE.scala 156:44 CSR.scala 19:23]
  wire [63:0] _GEN_136 = _is_mul_T ? mie : _GEN_129; // @[EXE.scala 156:44 CSR.scala 22:20]
  wire [63:0] _GEN_137 = _is_mul_T ? mip : _GEN_130; // @[EXE.scala 156:44 CSR.scala 23:20]
  wire [63:0] _GEN_138 = 7'h6d == io_in_bits_ctrl_signal_aluoptype ? _alu_result_T_7 : _GEN_131; // @[EXE.scala 156:44 179:18]
  wire [63:0] _GEN_139 = 7'h6d == io_in_bits_ctrl_signal_aluoptype ? mstatus : _GEN_132; // @[EXE.scala 156:44 CSR.scala 20:24]
  wire [63:0] _GEN_140 = 7'h6d == io_in_bits_ctrl_signal_aluoptype ? mtvec : _GEN_133; // @[EXE.scala 156:44 CSR.scala 21:22]
  wire [63:0] _GEN_141 = 7'h6d == io_in_bits_ctrl_signal_aluoptype ? mepc : _GEN_134; // @[EXE.scala 156:44 CSR.scala 18:17]
  wire [63:0] _GEN_142 = 7'h6d == io_in_bits_ctrl_signal_aluoptype ? mcause : _GEN_135; // @[EXE.scala 156:44 CSR.scala 19:23]
  wire [63:0] _GEN_143 = 7'h6d == io_in_bits_ctrl_signal_aluoptype ? mie : _GEN_136; // @[EXE.scala 156:44 CSR.scala 22:20]
  wire [63:0] _GEN_144 = 7'h6d == io_in_bits_ctrl_signal_aluoptype ? mip : _GEN_137; // @[EXE.scala 156:44 CSR.scala 23:20]
  wire [63:0] _GEN_145 = 7'h72 == io_in_bits_ctrl_signal_aluoptype ? _alu_result_T_12 : _GEN_138; // @[EXE.scala 156:44 176:18]
  wire [63:0] _GEN_146 = 7'h72 == io_in_bits_ctrl_signal_aluoptype ? mstatus : _GEN_139; // @[EXE.scala 156:44 CSR.scala 20:24]
  wire [63:0] _GEN_147 = 7'h72 == io_in_bits_ctrl_signal_aluoptype ? mtvec : _GEN_140; // @[EXE.scala 156:44 CSR.scala 21:22]
  wire [63:0] _GEN_148 = 7'h72 == io_in_bits_ctrl_signal_aluoptype ? mepc : _GEN_141; // @[EXE.scala 156:44 CSR.scala 18:17]
  wire [63:0] _GEN_149 = 7'h72 == io_in_bits_ctrl_signal_aluoptype ? mcause : _GEN_142; // @[EXE.scala 156:44 CSR.scala 19:23]
  wire [63:0] _GEN_150 = 7'h72 == io_in_bits_ctrl_signal_aluoptype ? mie : _GEN_143; // @[EXE.scala 156:44 CSR.scala 22:20]
  wire [63:0] _GEN_151 = 7'h72 == io_in_bits_ctrl_signal_aluoptype ? mip : _GEN_144; // @[EXE.scala 156:44 CSR.scala 23:20]
  wire [63:0] _GEN_152 = 7'h71 == io_in_bits_ctrl_signal_aluoptype ? _alu_result_T_11 : _GEN_145; // @[EXE.scala 156:44 173:18]
  wire [63:0] _GEN_153 = 7'h71 == io_in_bits_ctrl_signal_aluoptype ? mstatus : _GEN_146; // @[EXE.scala 156:44 CSR.scala 20:24]
  wire [63:0] _GEN_154 = 7'h71 == io_in_bits_ctrl_signal_aluoptype ? mtvec : _GEN_147; // @[EXE.scala 156:44 CSR.scala 21:22]
  wire [63:0] _GEN_155 = 7'h71 == io_in_bits_ctrl_signal_aluoptype ? mepc : _GEN_148; // @[EXE.scala 156:44 CSR.scala 18:17]
  wire [63:0] _GEN_156 = 7'h71 == io_in_bits_ctrl_signal_aluoptype ? mcause : _GEN_149; // @[EXE.scala 156:44 CSR.scala 19:23]
  wire [63:0] _GEN_157 = 7'h71 == io_in_bits_ctrl_signal_aluoptype ? mie : _GEN_150; // @[EXE.scala 156:44 CSR.scala 22:20]
  wire [63:0] _GEN_158 = 7'h71 == io_in_bits_ctrl_signal_aluoptype ? mip : _GEN_151; // @[EXE.scala 156:44 CSR.scala 23:20]
  wire [63:0] _GEN_159 = 7'h69 == io_in_bits_ctrl_signal_aluoptype ? _alu_result_T_10 : _GEN_152; // @[EXE.scala 156:44 170:18]
  wire [63:0] _GEN_160 = 7'h69 == io_in_bits_ctrl_signal_aluoptype ? mstatus : _GEN_153; // @[EXE.scala 156:44 CSR.scala 20:24]
  wire [63:0] _GEN_161 = 7'h69 == io_in_bits_ctrl_signal_aluoptype ? mtvec : _GEN_154; // @[EXE.scala 156:44 CSR.scala 21:22]
  wire [63:0] _GEN_162 = 7'h69 == io_in_bits_ctrl_signal_aluoptype ? mepc : _GEN_155; // @[EXE.scala 156:44 CSR.scala 18:17]
  wire [63:0] _GEN_163 = 7'h69 == io_in_bits_ctrl_signal_aluoptype ? mcause : _GEN_156; // @[EXE.scala 156:44 CSR.scala 19:23]
  wire [63:0] _GEN_164 = 7'h69 == io_in_bits_ctrl_signal_aluoptype ? mie : _GEN_157; // @[EXE.scala 156:44 CSR.scala 22:20]
  wire [63:0] _GEN_165 = 7'h69 == io_in_bits_ctrl_signal_aluoptype ? mip : _GEN_158; // @[EXE.scala 156:44 CSR.scala 23:20]
  wire [63:0] _GEN_166 = 7'h44 == io_in_bits_ctrl_signal_aluoptype ? _alu_result_T_8 : _GEN_159; // @[EXE.scala 156:44 167:18]
  wire [63:0] _GEN_167 = 7'h44 == io_in_bits_ctrl_signal_aluoptype ? mstatus : _GEN_160; // @[EXE.scala 156:44 CSR.scala 20:24]
  wire [63:0] _GEN_168 = 7'h44 == io_in_bits_ctrl_signal_aluoptype ? mtvec : _GEN_161; // @[EXE.scala 156:44 CSR.scala 21:22]
  wire [63:0] _GEN_169 = 7'h44 == io_in_bits_ctrl_signal_aluoptype ? mepc : _GEN_162; // @[EXE.scala 156:44 CSR.scala 18:17]
  wire [63:0] _GEN_170 = 7'h44 == io_in_bits_ctrl_signal_aluoptype ? mcause : _GEN_163; // @[EXE.scala 156:44 CSR.scala 19:23]
  wire [63:0] _GEN_171 = 7'h44 == io_in_bits_ctrl_signal_aluoptype ? mie : _GEN_164; // @[EXE.scala 156:44 CSR.scala 22:20]
  wire [63:0] _GEN_172 = 7'h44 == io_in_bits_ctrl_signal_aluoptype ? mip : _GEN_165; // @[EXE.scala 156:44 CSR.scala 23:20]
  wire [63:0] _GEN_173 = 7'h68 == io_in_bits_ctrl_signal_aluoptype ? _alu_result_T_7 : _GEN_166; // @[EXE.scala 156:44 164:18]
  wire [63:0] _GEN_174 = 7'h68 == io_in_bits_ctrl_signal_aluoptype ? mstatus : _GEN_167; // @[EXE.scala 156:44 CSR.scala 20:24]
  wire [63:0] _GEN_177 = 7'h68 == io_in_bits_ctrl_signal_aluoptype ? mcause : _GEN_170; // @[EXE.scala 156:44 CSR.scala 19:23]
  wire [63:0] _GEN_180 = 7'h1a == io_in_bits_ctrl_signal_aluoptype ? src2 : _GEN_173; // @[EXE.scala 156:44 161:18]
  wire [63:0] _GEN_181 = 7'h1a == io_in_bits_ctrl_signal_aluoptype ? mstatus : _GEN_174; // @[EXE.scala 156:44 CSR.scala 20:24]
  wire [63:0] alu_result = 7'h40 == io_in_bits_ctrl_signal_aluoptype ? _alu_result_T_1 : _GEN_180; // @[EXE.scala 156:44 158:18]
  wire [63:0] _shift_result_T = 3'h0 == io_in_bits_ctrl_signal_src1Type ? io_src1 : _GEN_1; // @[EXE.scala 226:29]
  wire [63:0] _shift_result_T_3 = $signed(_shift_result_T) >>> src2[4:0]; // @[EXE.scala 226:51]
  wire [94:0] _GEN_0 = {{31'd0}, src1}; // @[EXE.scala 230:39]
  wire [94:0] _shift_result_T_5 = _GEN_0 << src2[4:0]; // @[EXE.scala 230:39]
  wire  shift_result_sign = _shift_result_T_5[31]; // @[util.scala 11:19]
  wire [31:0] _shift_result_T_8 = shift_result_sign ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _shift_result_T_9 = {_shift_result_T_8,_shift_result_T_5[31:0]}; // @[Cat.scala 31:58]
  wire [126:0] _GEN_2 = {{63'd0}, src1}; // @[EXE.scala 233:28]
  wire [126:0] _shift_result_T_11 = _GEN_2 << src2[5:0]; // @[EXE.scala 233:28]
  wire [63:0] _shift_result_T_13 = src1 >> src2[5:0]; // @[EXE.scala 236:35]
  wire [94:0] _GEN_4 = {{63'd0}, src1[31:0]}; // @[EXE.scala 239:46]
  wire [94:0] _shift_result_T_16 = _GEN_4 << src2[5:0]; // @[EXE.scala 239:46]
  wire  shift_result_sign_1 = _shift_result_T_16[31]; // @[util.scala 11:19]
  wire [31:0] _shift_result_T_19 = shift_result_sign_1 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _shift_result_T_20 = {_shift_result_T_19,_shift_result_T_16[31:0]}; // @[Cat.scala 31:58]
  wire [31:0] _shift_result_T_22 = src1[31:0]; // @[EXE.scala 242:46]
  wire [31:0] _shift_result_T_25 = $signed(_shift_result_T_22) >>> src2[4:0]; // @[EXE.scala 242:68]
  wire  shift_result_sign_2 = _shift_result_T_25[31]; // @[util.scala 11:19]
  wire [31:0] _shift_result_T_27 = shift_result_sign_2 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _shift_result_T_28 = {_shift_result_T_27,_shift_result_T_25}; // @[Cat.scala 31:58]
  wire [31:0] _shift_result_T_31 = src1[31:0] >> src2[4:0]; // @[EXE.scala 245:46]
  wire  shift_result_sign_3 = _shift_result_T_31[31]; // @[util.scala 11:19]
  wire [31:0] _shift_result_T_34 = shift_result_sign_3 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _shift_result_T_35 = {_shift_result_T_34,_shift_result_T_31}; // @[Cat.scala 31:58]
  wire [63:0] _shift_result_T_54 = $signed(_shift_result_T) >>> src2[5:0]; // @[EXE.scala 254:51]
  wire [63:0] _GEN_194 = 7'h14 == io_in_bits_ctrl_signal_aluoptype ? _shift_result_T_54 : 64'h0; // @[EXE.scala 224:44 254:20]
  wire [63:0] _GEN_195 = 7'ha == io_in_bits_ctrl_signal_aluoptype ? _shift_result_T_35 : _GEN_194; // @[EXE.scala 224:44 251:20]
  wire [63:0] _GEN_196 = 7'h9 == io_in_bits_ctrl_signal_aluoptype ? _shift_result_T_28 : _GEN_195; // @[EXE.scala 224:44 248:20]
  wire [63:0] _GEN_197 = 7'h8 == io_in_bits_ctrl_signal_aluoptype ? _shift_result_T_35 : _GEN_196; // @[EXE.scala 224:44 245:20]
  wire [63:0] _GEN_198 = 7'h6 == io_in_bits_ctrl_signal_aluoptype ? _shift_result_T_28 : _GEN_197; // @[EXE.scala 224:44 242:20]
  wire [63:0] _GEN_199 = 7'h5 == io_in_bits_ctrl_signal_aluoptype ? _shift_result_T_20 : _GEN_198; // @[EXE.scala 224:44 239:20]
  wire [63:0] _GEN_200 = 7'h75 == io_in_bits_ctrl_signal_aluoptype ? _shift_result_T_13 : _GEN_199; // @[EXE.scala 224:44 236:20]
  wire [126:0] _GEN_201 = 7'h41 == io_in_bits_ctrl_signal_aluoptype ? _shift_result_T_11 : {{63'd0}, _GEN_200}; // @[EXE.scala 224:44 233:20]
  wire [126:0] _GEN_202 = 7'h73 == io_in_bits_ctrl_signal_aluoptype ? {{63'd0}, _shift_result_T_9} : _GEN_201; // @[EXE.scala 224:44 230:20]
  wire [126:0] _GEN_203 = 7'h6e == io_in_bits_ctrl_signal_aluoptype ? {{63'd0}, _shift_result_T_3} : _GEN_202; // @[EXE.scala 224:44 226:20]
  wire [63:0] _mul_io_in_bits_ctrl_data_src1_T_2 = {32'h0,src1[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _mul_io_in_bits_ctrl_data_src2_T_2 = {32'h0,src2[31:0]}; // @[Cat.scala 31:58]
  wire  _mul_io_in_valid_T = ~mul_io_out_valid; // @[EXE.scala 263:36]
  wire  div_io_in_bits_ctrl_data_src1_sign = src1[31]; // @[util.scala 11:19]
  wire [31:0] _div_io_in_bits_ctrl_data_src1_T_2 = div_io_in_bits_ctrl_data_src1_sign ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _div_io_in_bits_ctrl_data_src1_T_3 = {_div_io_in_bits_ctrl_data_src1_T_2,src1[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _div_io_in_bits_ctrl_data_src1_T_7 = is_div_sign ? _div_io_in_bits_ctrl_data_src1_T_3 :
    _mul_io_in_bits_ctrl_data_src1_T_2; // @[EXE.scala 269:51]
  wire  div_io_in_bits_ctrl_data_src2_sign = src2[31]; // @[util.scala 11:19]
  wire [31:0] _div_io_in_bits_ctrl_data_src2_T_2 = div_io_in_bits_ctrl_data_src2_sign ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _div_io_in_bits_ctrl_data_src2_T_3 = {_div_io_in_bits_ctrl_data_src2_T_2,src2[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _div_io_in_bits_ctrl_data_src2_T_7 = is_div_sign ? _div_io_in_bits_ctrl_data_src2_T_3 :
    _mul_io_in_bits_ctrl_data_src2_T_2; // @[EXE.scala 270:51]
  wire  _div_io_in_valid_T = ~div_io_out_valid; // @[EXE.scala 271:36]
  wire  _compar_result_T = src1 < src2; // @[EXE.scala 279:34]
  wire [63:0] _compar_result_T_1 = src1 < src2 ? 64'h1 : 64'h0; // @[EXE.scala 279:27]
  wire [63:0] _compar_result_T_3 = 3'h0 == io_in_bits_ctrl_signal_src2Type ? io_src2 : _GEN_3; // @[EXE.scala 282:48]
  wire  _compar_result_T_4 = $signed(_shift_result_T) < $signed(_compar_result_T_3); // @[EXE.scala 282:41]
  wire [63:0] _compar_result_T_5 = $signed(_shift_result_T) < $signed(_compar_result_T_3) ? 64'h1 : 64'h0; // @[EXE.scala 282:27]
  wire [63:0] _GEN_204 = 7'h2 == io_in_bits_ctrl_signal_aluoptype ? _compar_result_T_5 : 64'h0; // @[EXE.scala 277:44 282:21]
  wire [63:0] compar_result = 7'h6a == io_in_bits_ctrl_signal_aluoptype ? _compar_result_T_1 : _GEN_204; // @[EXE.scala 277:44 279:21]
  wire  _jump_result_T = io_in_bits_ctrl_signal_fuType == 3'h3; // @[EXE.scala 287:52]
  wire [63:0] jump_result = io_in_bits_ctrl_signal_fuType == 3'h3 ? _dnpc_T_1 : 64'h0; // @[EXE.scala 287:21]
  wire [63:0] _GEN_206 = 3'h5 == io_in_bits_ctrl_signal_fuType ? compar_result : 64'h0; // @[EXE.scala 290:41 304:18]
  wire [63:0] shift_result = _GEN_203[63:0];
  wire [63:0] _GEN_207 = 3'h1 == io_in_bits_ctrl_signal_fuType ? shift_result : _GEN_206; // @[EXE.scala 290:41 301:18]
  wire [63:0] _GEN_208 = 3'h2 == io_in_bits_ctrl_signal_fuType ? 64'h0 : _GEN_207; // @[EXE.scala 290:41 298:18]
  wire [63:0] _GEN_209 = 3'h3 == io_in_bits_ctrl_signal_fuType ? jump_result : _GEN_208; // @[EXE.scala 290:41 295:18]
  wire  _T_71 = 7'h6b == io_in_bits_ctrl_signal_aluoptype; // @[EXE.scala 312:44]
  wire [63:0] _branch_result_T_1 = io_in_bits_ctrl_flow_PC + io_in_bits_ctrl_data_Imm; // @[EXE.scala 314:27]
  wire  _T_72 = 7'h6c == io_in_bits_ctrl_signal_aluoptype; // @[EXE.scala 312:44]
  wire  _T_73 = 7'h76 == io_in_bits_ctrl_signal_aluoptype; // @[EXE.scala 312:44]
  wire  _T_74 = 7'h7b == io_in_bits_ctrl_signal_aluoptype; // @[EXE.scala 312:44]
  wire  _T_75 = 7'hb == io_in_bits_ctrl_signal_aluoptype; // @[EXE.scala 312:44]
  wire  _T_76 = 7'hc == io_in_bits_ctrl_signal_aluoptype; // @[EXE.scala 312:44]
  wire  _T_77 = 7'h17 == io_in_bits_ctrl_signal_aluoptype; // @[EXE.scala 312:44]
  wire  _T_78 = 7'h18 == io_in_bits_ctrl_signal_aluoptype; // @[EXE.scala 312:44]
  wire  _GEN_212 = 7'h17 == io_in_bits_ctrl_signal_aluoptype | 7'h18 == io_in_bits_ctrl_signal_aluoptype; // @[EXE.scala 312:44 339:19]
  wire [63:0] _GEN_213 = 7'hc == io_in_bits_ctrl_signal_aluoptype ? _branch_result_T_1 : 64'h0; // @[EXE.scala 312:44 334:21]
  wire  _GEN_214 = 7'hc == io_in_bits_ctrl_signal_aluoptype ? src1 >= src2 : _GEN_212; // @[EXE.scala 312:44 335:19]
  wire [63:0] _GEN_215 = 7'hb == io_in_bits_ctrl_signal_aluoptype ? _branch_result_T_1 : _GEN_213; // @[EXE.scala 312:44 330:21]
  wire  _GEN_216 = 7'hb == io_in_bits_ctrl_signal_aluoptype ? _compar_result_T : _GEN_214; // @[EXE.scala 312:44 331:19]
  wire [63:0] _GEN_217 = 7'h7b == io_in_bits_ctrl_signal_aluoptype ? _branch_result_T_1 : _GEN_215; // @[EXE.scala 312:44 326:21]
  wire  _GEN_218 = 7'h7b == io_in_bits_ctrl_signal_aluoptype ? _compar_result_T_4 : _GEN_216; // @[EXE.scala 312:44 327:19]
  wire [63:0] _GEN_219 = 7'h76 == io_in_bits_ctrl_signal_aluoptype ? _branch_result_T_1 : _GEN_217; // @[EXE.scala 312:44 322:21]
  wire  _GEN_220 = 7'h76 == io_in_bits_ctrl_signal_aluoptype ? $signed(_shift_result_T) >= $signed(_compar_result_T_3)
     : _GEN_218; // @[EXE.scala 312:44 323:19]
  wire [63:0] _GEN_221 = 7'h6c == io_in_bits_ctrl_signal_aluoptype ? _branch_result_T_1 : _GEN_219; // @[EXE.scala 312:44 318:21]
  wire  _GEN_222 = 7'h6c == io_in_bits_ctrl_signal_aluoptype ? src1 != src2 : _GEN_220; // @[EXE.scala 312:44 319:19]
  wire [63:0] branch_result = 7'h6b == io_in_bits_ctrl_signal_aluoptype ? _branch_result_T_1 : _GEN_221; // @[EXE.scala 312:44 314:21]
  wire  branch_flag = 7'h6b == io_in_bits_ctrl_signal_aluoptype ? src1 == src2 : _GEN_222; // @[EXE.scala 312:44 315:19]
  wire [63:0] _T_92 = mstatus & 64'hfffffffffffffff7; // @[EXE.scala 350:64]
  wire [63:0] _T_112 = mstatus | 64'h8; // @[EXE.scala 354:64]
  wire [63:0] _GEN_267 = _T_78 ? mepc : 64'h0; // @[EXE.scala 347:44 353:16]
  wire [63:0] csr_data = _T_77 ? mtvec : _GEN_267; // @[EXE.scala 347:44 349:16]
  wire [63:0] _dnpc_T_7 = {_alu_result_T_1[63:1],1'h0}; // @[Cat.scala 31:58]
  wire [63:0] _dnpc_T_11 = branch_flag ? branch_result : _dnpc_T_1; // @[EXE.scala 367:18]
  wire [63:0] _GEN_281 = _T_78 ? csr_data : _dnpc_T_1; // @[EXE.scala 359:44 390:12]
  wire [63:0] _GEN_282 = _T_77 ? csr_data : _GEN_281; // @[EXE.scala 359:44 387:12]
  wire [63:0] _GEN_283 = _T_75 ? _dnpc_T_11 : _GEN_282; // @[EXE.scala 359:44 383:12]
  wire [63:0] _GEN_284 = _T_74 ? _dnpc_T_11 : _GEN_283; // @[EXE.scala 359:44 380:12]
  wire [63:0] _GEN_285 = _T_76 ? _dnpc_T_11 : _GEN_284; // @[EXE.scala 359:44 377:12]
  wire [63:0] _GEN_286 = _T_73 ? _dnpc_T_11 : _GEN_285; // @[EXE.scala 359:44 374:12]
  wire [63:0] _GEN_287 = _T_72 ? _dnpc_T_11 : _GEN_286; // @[EXE.scala 359:44 371:12]
  wire [63:0] _GEN_288 = _T_71 ? _dnpc_T_11 : _GEN_287; // @[EXE.scala 359:44 367:12]
  wire [63:0] _GEN_289 = 7'h48 == io_in_bits_ctrl_signal_aluoptype ? _dnpc_T_7 : _GEN_288; // @[EXE.scala 359:44 364:12]
  reg [63:0] CSRDIFF_io_mtvec_REG; // @[EXE.scala 409:38]
  reg [63:0] CSRDIFF_io_mtvec_REG_1; // @[EXE.scala 409:30]
  reg [63:0] CSRDIFF_io_mcause_REG; // @[EXE.scala 410:39]
  reg [63:0] CSRDIFF_io_mcause_REG_1; // @[EXE.scala 410:31]
  reg [63:0] CSRDIFF_io_mepc_REG; // @[EXE.scala 411:37]
  reg [63:0] CSRDIFF_io_mepc_REG_1; // @[EXE.scala 411:29]
  reg [63:0] CSRDIFF_io_mstatus_REG; // @[EXE.scala 412:40]
  reg [63:0] CSRDIFF_io_mstatus_REG_1; // @[EXE.scala 412:32]
  wire  _io_out_valid_T_1 = _mul_io_in_valid_T & is_mul; // @[EXE.scala 436:43]
  wire  _io_out_valid_T_4 = _div_io_in_valid_T & is_div; // @[EXE.scala 436:78]
  CSR_DIFF CSRDIFF ( // @[EXE.scala 115:21]
    .mepc(CSRDIFF_mepc),
    .mcause(CSRDIFF_mcause),
    .mstatus(CSRDIFF_mstatus),
    .mtvec(CSRDIFF_mtvec)
  );
  MUL mul ( // @[EXE.scala 118:19]
    .clock(mul_clock),
    .reset(mul_reset),
    .io_in_valid(mul_io_in_valid),
    .io_in_bits_ctrl_data_src1(mul_io_in_bits_ctrl_data_src1),
    .io_in_bits_ctrl_data_src2(mul_io_in_bits_ctrl_data_src2),
    .io_out_valid(mul_io_out_valid),
    .io_out_bits_result_result_lo(mul_io_out_bits_result_result_lo)
  );
  DIV div ( // @[EXE.scala 119:19]
    .clock(div_clock),
    .reset(div_reset),
    .io_in_valid(div_io_in_valid),
    .io_in_bits_ctrl_flow_div_signed(div_io_in_bits_ctrl_flow_div_signed),
    .io_in_bits_ctrl_data_src1(div_io_in_bits_ctrl_data_src1),
    .io_in_bits_ctrl_data_src2(div_io_in_bits_ctrl_data_src2),
    .io_out_valid(div_io_out_valid),
    .io_out_bits_result_quotient(div_io_out_bits_result_quotient),
    .io_out_bits_result_remainder(div_io_out_bits_result_remainder)
  );
  assign io_in_ready = (_io_out_valid_T_1 | _io_out_valid_T_4) & io_in_valid ? 1'h0 : io_out_ready; // @[EXE.scala 437:21]
  assign io_branchIO_is_branch = branch_flag & io_out_bits_ctrl_signal_inst_valid & io_in_valid & io_out_ready; // @[EXE.scala 433:91]
  assign io_branchIO_is_jump = _jump_result_T & io_out_bits_ctrl_signal_inst_valid & io_in_valid & io_out_ready; // @[EXE.scala 434:129]
  assign io_branchIO_dnpc = 7'h19 == io_in_bits_ctrl_signal_aluoptype ? _alu_result_T_1 : _GEN_289; // @[EXE.scala 359:44 361:12]
  assign io_out_valid = ~(_mul_io_in_valid_T & is_mul) & ~(_div_io_in_valid_T & is_div) & io_in_valid; // @[EXE.scala 436:89]
  assign io_out_bits_ctrl_signal_fuType = io_in_bits_ctrl_signal_fuType; // @[EXE.scala 419:27]
  assign io_out_bits_ctrl_signal_inst_valid = io_in_bits_ctrl_signal_inst_valid; // @[EXE.scala 423:38]
  assign io_out_bits_ctrl_signal_rfWen = io_in_bits_ctrl_signal_rfWen; // @[EXE.scala 419:27]
  assign io_out_bits_ctrl_signal_aluoptype = io_in_bits_ctrl_signal_aluoptype; // @[EXE.scala 419:27]
  assign io_out_bits_ctrl_flow_PC = io_in_bits_ctrl_flow_PC; // @[EXE.scala 420:25]
  assign io_out_bits_ctrl_flow_inst = io_in_bits_ctrl_flow_inst; // @[EXE.scala 420:25]
  assign io_out_bits_ctrl_flow_Dnpc = 7'h19 == io_in_bits_ctrl_signal_aluoptype ? _alu_result_T_1 : _GEN_289; // @[EXE.scala 359:44 361:12]
  assign io_out_bits_ctrl_rf_rfDest = io_in_bits_ctrl_signal_rfDest; // @[EXE.scala 429:30]
  assign io_out_bits_ctrl_rf_rfWen = io_in_valid & io_in_bits_ctrl_signal_rfWen; // @[EXE.scala 430:35]
  assign io_out_bits_ctrl_rf_rfData = 3'h0 == io_in_bits_ctrl_signal_fuType ? alu_result : _GEN_209; // @[EXE.scala 290:41 292:18]
  assign io_out_bits_ctrl_data_src1 = 3'h0 == io_in_bits_ctrl_signal_src1Type ? io_src1 : _GEN_1; // @[EXE.scala 124:43 126:12]
  assign io_out_bits_ctrl_data_src2 = 3'h0 == io_in_bits_ctrl_signal_src2Type ? io_src2 : _GEN_3; // @[EXE.scala 135:43 138:12]
  assign io_out_bits_ctrl_data_Imm = io_in_bits_ctrl_data_Imm; // @[EXE.scala 421:25]
  assign io_is_break = io_in_bits_ctrl_signal_aluoptype == 7'h42 & io_out_bits_ctrl_signal_inst_valid; // @[EXE.scala 415:77]
  assign io_is_flush = (branch_flag | io_branchIO_is_jump) & io_in_valid; // @[EXE.scala 414:75]
  assign CSRDIFF_mepc = CSRDIFF_io_mepc_REG_1; // @[EXE.scala 411:19]
  assign CSRDIFF_mcause = CSRDIFF_io_mcause_REG_1; // @[EXE.scala 410:21]
  assign CSRDIFF_mstatus = CSRDIFF_io_mstatus_REG_1; // @[EXE.scala 412:22]
  assign CSRDIFF_mtvec = CSRDIFF_io_mtvec_REG_1; // @[EXE.scala 409:20]
  assign mul_clock = clock;
  assign mul_reset = reset;
  assign mul_io_in_valid = is_mul & ~mul_io_out_valid; // @[EXE.scala 263:33]
  assign mul_io_in_bits_ctrl_data_src1 = is_mul ? src1 : _mul_io_in_bits_ctrl_data_src1_T_2; // @[EXE.scala 259:39]
  assign mul_io_in_bits_ctrl_data_src2 = is_mul ? src2 : _mul_io_in_bits_ctrl_data_src2_T_2; // @[EXE.scala 260:39]
  assign div_clock = clock;
  assign div_reset = reset;
  assign div_io_in_valid = is_div & ~div_io_out_valid; // @[EXE.scala 271:33]
  assign div_io_in_bits_ctrl_flow_div_signed = _is_div_sign_T_2 | _is_div_T_7 | _is_div_T_11; // @[EXE.scala 112:59]
  assign div_io_in_bits_ctrl_data_src1 = is_divw ? _div_io_in_bits_ctrl_data_src1_T_7 : src1; // @[EXE.scala 269:39]
  assign div_io_in_bits_ctrl_data_src2 = is_divw ? _div_io_in_bits_ctrl_data_src2_T_7 : src2; // @[EXE.scala 270:39]
  always @(posedge clock) begin
    if (_T_77) begin // @[EXE.scala 394:44]
      mepc <= io_in_bits_ctrl_flow_PC;
    end else if (!(7'h40 == io_in_bits_ctrl_signal_aluoptype)) begin // @[EXE.scala 156:44]
      if (!(7'h1a == io_in_bits_ctrl_signal_aluoptype)) begin // @[EXE.scala 156:44]
        if (!(7'h68 == io_in_bits_ctrl_signal_aluoptype)) begin // @[EXE.scala 156:44]
          mepc <= _GEN_169;
        end
      end
    end
    if (reset) begin // @[CSR.scala 19:23]
      mcause <= 64'h0; // @[CSR.scala 19:23]
    end else if (_T_77) begin // @[EXE.scala 394:44]
      mcause <= 64'hb;
    end else if (!(7'h40 == io_in_bits_ctrl_signal_aluoptype)) begin // @[EXE.scala 156:44]
      if (!(7'h1a == io_in_bits_ctrl_signal_aluoptype)) begin // @[EXE.scala 156:44]
        mcause <= _GEN_177;
      end
    end
    if (reset) begin // @[CSR.scala 20:24]
      mstatus <= 64'h0; // @[CSR.scala 20:24]
    end else if (_T_77) begin // @[EXE.scala 347:44]
      mstatus <= _T_92;
    end else if (_T_78) begin // @[EXE.scala 347:44]
      mstatus <= _T_112;
    end else if (!(7'h40 == io_in_bits_ctrl_signal_aluoptype)) begin // @[EXE.scala 156:44]
      mstatus <= _GEN_181;
    end
    if (reset) begin // @[CSR.scala 21:22]
      mtvec <= 64'h0; // @[CSR.scala 21:22]
    end else if (!(7'h40 == io_in_bits_ctrl_signal_aluoptype)) begin // @[EXE.scala 156:44]
      if (!(7'h1a == io_in_bits_ctrl_signal_aluoptype)) begin // @[EXE.scala 156:44]
        if (!(7'h68 == io_in_bits_ctrl_signal_aluoptype)) begin // @[EXE.scala 156:44]
          mtvec <= _GEN_168;
        end
      end
    end
    if (reset) begin // @[CSR.scala 22:20]
      mie <= 64'h0; // @[CSR.scala 22:20]
    end else if (!(7'h40 == io_in_bits_ctrl_signal_aluoptype)) begin // @[EXE.scala 156:44]
      if (!(7'h1a == io_in_bits_ctrl_signal_aluoptype)) begin // @[EXE.scala 156:44]
        if (!(7'h68 == io_in_bits_ctrl_signal_aluoptype)) begin // @[EXE.scala 156:44]
          mie <= _GEN_171;
        end
      end
    end
    if (reset) begin // @[CSR.scala 23:20]
      mip <= 64'h0; // @[CSR.scala 23:20]
    end else if (!(7'h40 == io_in_bits_ctrl_signal_aluoptype)) begin // @[EXE.scala 156:44]
      if (!(7'h1a == io_in_bits_ctrl_signal_aluoptype)) begin // @[EXE.scala 156:44]
        if (!(7'h68 == io_in_bits_ctrl_signal_aluoptype)) begin // @[EXE.scala 156:44]
          mip <= _GEN_172;
        end
      end
    end
    CSRDIFF_io_mtvec_REG <= mtvec; // @[EXE.scala 409:38]
    CSRDIFF_io_mtvec_REG_1 <= CSRDIFF_io_mtvec_REG; // @[EXE.scala 409:30]
    CSRDIFF_io_mcause_REG <= mcause; // @[EXE.scala 410:39]
    CSRDIFF_io_mcause_REG_1 <= CSRDIFF_io_mcause_REG; // @[EXE.scala 410:31]
    CSRDIFF_io_mepc_REG <= mepc; // @[EXE.scala 411:37]
    CSRDIFF_io_mepc_REG_1 <= CSRDIFF_io_mepc_REG; // @[EXE.scala 411:29]
    CSRDIFF_io_mstatus_REG <= mstatus; // @[EXE.scala 412:40]
    CSRDIFF_io_mstatus_REG_1 <= CSRDIFF_io_mstatus_REG; // @[EXE.scala 412:32]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mepc = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mcause = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mstatus = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mtvec = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mie = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mip = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  CSRDIFF_io_mtvec_REG = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  CSRDIFF_io_mtvec_REG_1 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  CSRDIFF_io_mcause_REG = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  CSRDIFF_io_mcause_REG_1 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  CSRDIFF_io_mepc_REG = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  CSRDIFF_io_mepc_REG_1 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  CSRDIFF_io_mstatus_REG = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  CSRDIFF_io_mstatus_REG_1 = _RAND_13[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MEM_stage(
  output        io_in_ready,
  input         io_in_valid,
  input  [2:0]  io_in_bits_ctrl_signal_fuType,
  input         io_in_bits_ctrl_signal_inst_valid,
  input         io_in_bits_ctrl_signal_rfWen,
  input  [6:0]  io_in_bits_ctrl_signal_aluoptype,
  input  [63:0] io_in_bits_ctrl_flow_PC,
  input  [31:0] io_in_bits_ctrl_flow_inst,
  input  [63:0] io_in_bits_ctrl_flow_Dnpc,
  input  [4:0]  io_in_bits_ctrl_rf_rfDest,
  input  [63:0] io_in_bits_ctrl_rf_rfData,
  input  [63:0] io_in_bits_ctrl_data_src1,
  input  [63:0] io_in_bits_ctrl_data_src2,
  input  [63:0] io_in_bits_ctrl_data_Imm,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_ctrl_signal_inst_valid,
  output        io_out_bits_ctrl_signal_rfWen,
  output [63:0] io_out_bits_ctrl_flow_PC,
  output [31:0] io_out_bits_ctrl_flow_inst,
  output [63:0] io_out_bits_ctrl_flow_Dnpc,
  output        io_out_bits_ctrl_flow_skip,
  output [4:0]  io_out_bits_ctrl_rf_rfDest,
  output        io_out_bits_ctrl_rf_rfWen,
  output [63:0] io_out_bits_ctrl_rf_rfData,
  output        io_cache_io_addr_req_valid,
  output [63:0] io_cache_io_addr_req_bits_addr,
  output        io_cache_io_addr_req_bits_ce,
  output        io_cache_io_addr_req_bits_we,
  input         io_cache_io_rdata_rep_valid,
  input  [63:0] io_cache_io_rdata_rep_bits_rdata,
  output [63:0] io_cache_io_wdata_req_bits_wdata,
  output [7:0]  io_cache_io_wdata_req_bits_wmask,
  input         io_cache_io_wdata_rep
);
  wire  _T_62 = 7'h45 == io_in_bits_ctrl_signal_aluoptype; // @[MEM.scala 54:44]
  wire [63:0] _addr_temp_T_1 = io_in_bits_ctrl_data_src1 + io_in_bits_ctrl_data_Imm; // @[MEM.scala 56:25]
  wire  _T_63 = 7'h46 == io_in_bits_ctrl_signal_aluoptype; // @[MEM.scala 54:44]
  wire  _T_64 = 7'h70 == io_in_bits_ctrl_signal_aluoptype; // @[MEM.scala 54:44]
  wire  _T_65 = 7'h47 == io_in_bits_ctrl_signal_aluoptype; // @[MEM.scala 54:44]
  wire  _T_66 = 7'h11 == io_in_bits_ctrl_signal_aluoptype; // @[MEM.scala 54:44]
  wire  _T_67 = 7'h6f == io_in_bits_ctrl_signal_aluoptype; // @[MEM.scala 54:44]
  wire  _T_68 = 7'he == io_in_bits_ctrl_signal_aluoptype; // @[MEM.scala 54:44]
  wire  _T_69 = 7'h74 == io_in_bits_ctrl_signal_aluoptype; // @[MEM.scala 54:44]
  wire  _T_70 = 7'h77 == io_in_bits_ctrl_signal_aluoptype; // @[MEM.scala 54:44]
  wire  _T_71 = 7'h3 == io_in_bits_ctrl_signal_aluoptype; // @[MEM.scala 54:44]
  wire  _T_72 = 7'h4 == io_in_bits_ctrl_signal_aluoptype; // @[MEM.scala 54:44]
  wire [63:0] _GEN_0 = 7'h4 == io_in_bits_ctrl_signal_aluoptype ? _addr_temp_T_1 : 64'h0; // @[MEM.scala 54:44 90:17]
  wire [63:0] _GEN_1 = 7'h3 == io_in_bits_ctrl_signal_aluoptype ? _addr_temp_T_1 : _GEN_0; // @[MEM.scala 54:44 87:17]
  wire [63:0] _GEN_2 = 7'h77 == io_in_bits_ctrl_signal_aluoptype ? _addr_temp_T_1 : _GEN_1; // @[MEM.scala 54:44 83:17]
  wire [63:0] _GEN_4 = 7'h74 == io_in_bits_ctrl_signal_aluoptype ? _addr_temp_T_1 : _GEN_2; // @[MEM.scala 54:44 79:17]
  wire [63:0] _GEN_6 = 7'he == io_in_bits_ctrl_signal_aluoptype ? _addr_temp_T_1 : _GEN_4; // @[MEM.scala 54:44 76:17]
  wire [63:0] _GEN_8 = 7'h6f == io_in_bits_ctrl_signal_aluoptype ? _addr_temp_T_1 : _GEN_6; // @[MEM.scala 54:44 73:17]
  wire [63:0] _GEN_10 = 7'h11 == io_in_bits_ctrl_signal_aluoptype ? _addr_temp_T_1 : _GEN_8; // @[MEM.scala 54:44 70:17]
  wire [63:0] _GEN_12 = 7'h47 == io_in_bits_ctrl_signal_aluoptype ? _addr_temp_T_1 : _GEN_10; // @[MEM.scala 54:44 67:17]
  wire [63:0] _GEN_14 = 7'h70 == io_in_bits_ctrl_signal_aluoptype ? _addr_temp_T_1 : _GEN_12; // @[MEM.scala 54:44 63:17]
  wire [63:0] _GEN_16 = 7'h46 == io_in_bits_ctrl_signal_aluoptype ? _addr_temp_T_1 : _GEN_14; // @[MEM.scala 54:44 59:17]
  wire [63:0] addr_temp = 7'h45 == io_in_bits_ctrl_signal_aluoptype ? _addr_temp_T_1 : _GEN_16; // @[MEM.scala 54:44 56:17]
  wire  _T_1 = addr_temp[2:0] == 3'h0; // @[MEM.scala 34:22]
  wire  _T_3 = addr_temp[2:0] == 3'h1; // @[MEM.scala 35:22]
  wire  _T_5 = addr_temp[2:0] == 3'h2; // @[MEM.scala 36:22]
  wire  _T_7 = addr_temp[2:0] == 3'h3; // @[MEM.scala 37:22]
  wire  _T_9 = addr_temp[2:0] == 3'h4; // @[MEM.scala 38:22]
  wire  _T_11 = addr_temp[2:0] == 3'h5; // @[MEM.scala 39:22]
  wire  _T_13 = addr_temp[2:0] == 3'h6; // @[MEM.scala 40:22]
  wire  _T_15 = addr_temp[2:0] == 3'h7; // @[MEM.scala 41:22]
  wire [63:0] _T_20 = {56'h0,io_in_bits_ctrl_data_src2[7:0]}; // @[Cat.scala 31:58]
  wire [63:0] _T_26 = {48'h0,io_in_bits_ctrl_data_src2[7:0],8'h0}; // @[Cat.scala 31:58]
  wire [63:0] _T_32 = {40'h0,io_in_bits_ctrl_data_src2[7:0],16'h0}; // @[Cat.scala 31:58]
  wire [63:0] _T_38 = {32'h0,io_in_bits_ctrl_data_src2[7:0],24'h0}; // @[Cat.scala 31:58]
  wire [63:0] _T_44 = {24'h0,io_in_bits_ctrl_data_src2[7:0],32'h0}; // @[Cat.scala 31:58]
  wire [63:0] _T_50 = {16'h0,io_in_bits_ctrl_data_src2[7:0],40'h0}; // @[Cat.scala 31:58]
  wire [63:0] _T_56 = {8'h0,io_in_bits_ctrl_data_src2[7:0],48'h0}; // @[Cat.scala 31:58]
  wire [63:0] _T_61 = {io_in_bits_ctrl_data_src2[7:0],56'h0}; // @[Cat.scala 31:58]
  wire  _GEN_5 = 7'h74 == io_in_bits_ctrl_signal_aluoptype | 7'h77 == io_in_bits_ctrl_signal_aluoptype; // @[MEM.scala 54:44 80:10]
  wire  _GEN_7 = 7'he == io_in_bits_ctrl_signal_aluoptype ? 1'h0 : _GEN_5; // @[MEM.scala 54:44]
  wire  _GEN_9 = 7'h6f == io_in_bits_ctrl_signal_aluoptype ? 1'h0 : _GEN_7; // @[MEM.scala 54:44]
  wire  _GEN_11 = 7'h11 == io_in_bits_ctrl_signal_aluoptype ? 1'h0 : _GEN_9; // @[MEM.scala 54:44]
  wire  _GEN_13 = 7'h47 == io_in_bits_ctrl_signal_aluoptype ? 1'h0 : _GEN_11; // @[MEM.scala 54:44]
  wire  _GEN_15 = 7'h70 == io_in_bits_ctrl_signal_aluoptype | _GEN_13; // @[MEM.scala 54:44 64:10]
  wire  _GEN_17 = 7'h46 == io_in_bits_ctrl_signal_aluoptype | _GEN_15; // @[MEM.scala 54:44 60:10]
  wire [63:0] _wdata_temp_T_2 = {48'h0,io_in_bits_ctrl_data_src2[15:0]}; // @[Cat.scala 31:58]
  wire [63:0] _wdata_temp_T_6 = {32'h0,io_in_bits_ctrl_data_src2[15:0],16'h0}; // @[Cat.scala 31:58]
  wire [63:0] _wdata_temp_T_10 = {16'h0,io_in_bits_ctrl_data_src2[15:0],32'h0}; // @[Cat.scala 31:58]
  wire [63:0] _wdata_temp_T_13 = {io_in_bits_ctrl_data_src2[15:0],48'h0}; // @[Cat.scala 31:58]
  wire [7:0] _GEN_20 = 2'h3 == addr_temp[2:1] ? 8'hc0 : 8'h0; // @[MEM.scala 100:31 114:22]
  wire [63:0] _GEN_21 = 2'h3 == addr_temp[2:1] ? _wdata_temp_T_13 : 64'h0; // @[MEM.scala 100:31 115:22]
  wire [7:0] _GEN_22 = 2'h2 == addr_temp[2:1] ? 8'h30 : _GEN_20; // @[MEM.scala 100:31 110:22]
  wire [63:0] _GEN_23 = 2'h2 == addr_temp[2:1] ? _wdata_temp_T_10 : _GEN_21; // @[MEM.scala 100:31 111:22]
  wire [7:0] _GEN_24 = 2'h1 == addr_temp[2:1] ? 8'hc : _GEN_22; // @[MEM.scala 100:31 106:22]
  wire [63:0] _GEN_25 = 2'h1 == addr_temp[2:1] ? _wdata_temp_T_6 : _GEN_23; // @[MEM.scala 100:31 107:22]
  wire [7:0] _GEN_26 = 2'h0 == addr_temp[2:1] ? 8'h3 : _GEN_24; // @[MEM.scala 100:31 102:22]
  wire [63:0] _GEN_27 = 2'h0 == addr_temp[2:1] ? _wdata_temp_T_2 : _GEN_25; // @[MEM.scala 100:31 103:22]
  wire [7:0] _wmask_temp_T = _T_15 ? 8'h80 : 8'h0; // @[Mux.scala 101:16]
  wire [7:0] _wmask_temp_T_1 = _T_13 ? 8'h40 : _wmask_temp_T; // @[Mux.scala 101:16]
  wire [7:0] _wmask_temp_T_2 = _T_11 ? 8'h20 : _wmask_temp_T_1; // @[Mux.scala 101:16]
  wire [7:0] _wmask_temp_T_3 = _T_9 ? 8'h10 : _wmask_temp_T_2; // @[Mux.scala 101:16]
  wire [7:0] _wmask_temp_T_4 = _T_7 ? 8'h8 : _wmask_temp_T_3; // @[Mux.scala 101:16]
  wire [7:0] _wmask_temp_T_5 = _T_5 ? 8'h4 : _wmask_temp_T_4; // @[Mux.scala 101:16]
  wire [7:0] _wmask_temp_T_6 = _T_3 ? 8'h2 : _wmask_temp_T_5; // @[Mux.scala 101:16]
  wire [7:0] _wmask_temp_T_7 = _T_1 ? 8'h1 : _wmask_temp_T_6; // @[Mux.scala 101:16]
  wire [63:0] _wdata_temp_T_14 = _T_15 ? _T_61 : 64'h0; // @[Mux.scala 101:16]
  wire [63:0] _wdata_temp_T_15 = _T_13 ? _T_56 : _wdata_temp_T_14; // @[Mux.scala 101:16]
  wire [63:0] _wdata_temp_T_16 = _T_11 ? _T_50 : _wdata_temp_T_15; // @[Mux.scala 101:16]
  wire [63:0] _wdata_temp_T_17 = _T_9 ? _T_44 : _wdata_temp_T_16; // @[Mux.scala 101:16]
  wire [63:0] _wdata_temp_T_18 = _T_7 ? _T_38 : _wdata_temp_T_17; // @[Mux.scala 101:16]
  wire [63:0] _wdata_temp_T_19 = _T_5 ? _T_32 : _wdata_temp_T_18; // @[Mux.scala 101:16]
  wire [63:0] _wdata_temp_T_20 = _T_3 ? _T_26 : _wdata_temp_T_19; // @[Mux.scala 101:16]
  wire [63:0] _wdata_temp_T_21 = _T_1 ? _T_20 : _wdata_temp_T_20; // @[Mux.scala 101:16]
  wire [7:0] _wmask_temp_T_10 = addr_temp[2] ? 8'hf0 : 8'hf; // @[MEM.scala 125:24]
  wire [63:0] _wdata_temp_T_26 = {io_in_bits_ctrl_data_src2[31:0],32'h0}; // @[Cat.scala 31:58]
  wire [63:0] _wdata_temp_T_29 = {32'h0,io_in_bits_ctrl_data_src2[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _wdata_temp_T_30 = addr_temp[2] ? _wdata_temp_T_26 : _wdata_temp_T_29; // @[MEM.scala 126:24]
  wire [7:0] _GEN_28 = _T_70 ? _wmask_temp_T_10 : 8'h0; // @[MEM.scala 125:18 93:44]
  wire [63:0] _GEN_29 = _T_70 ? _wdata_temp_T_30 : 64'h0; // @[MEM.scala 126:18 93:44]
  wire [7:0] _GEN_30 = _T_69 ? _wmask_temp_T_7 : _GEN_28; // @[MEM.scala 121:18 93:44]
  wire [63:0] _GEN_31 = _T_69 ? _wdata_temp_T_21 : _GEN_29; // @[MEM.scala 122:18 93:44]
  wire [7:0] _GEN_32 = _T_64 ? _GEN_26 : _GEN_30; // @[MEM.scala 93:44]
  wire [63:0] _GEN_33 = _T_64 ? _GEN_27 : _GEN_31; // @[MEM.scala 93:44]
  wire  _T_107 = addr_temp[2:1] == 2'h0; // @[MEM.scala 140:22]
  wire  _T_110 = addr_temp[2:1] == 2'h1; // @[MEM.scala 141:22]
  wire  _T_113 = addr_temp[2:1] == 2'h2; // @[MEM.scala 142:22]
  wire  _T_116 = addr_temp[2:1] == 2'h3; // @[MEM.scala 143:22]
  wire  mem_result_sign = io_cache_io_rdata_rep_bits_rdata[63]; // @[util.scala 11:19]
  wire [31:0] _mem_result_T_4 = mem_result_sign ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _mem_result_T_5 = {_mem_result_T_4,io_cache_io_rdata_rep_bits_rdata[63:32]}; // @[Cat.scala 31:58]
  wire  mem_result_sign_1 = io_cache_io_rdata_rep_bits_rdata[31]; // @[util.scala 11:19]
  wire [31:0] _mem_result_T_8 = mem_result_sign_1 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _mem_result_T_9 = {_mem_result_T_8,io_cache_io_rdata_rep_bits_rdata[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _mem_result_T_10 = addr_temp[2] ? _mem_result_T_5 : _mem_result_T_9; // @[MEM.scala 151:24]
  wire [63:0] _mem_result_T_15 = {32'h0,io_cache_io_rdata_rep_bits_rdata[63:32]}; // @[Cat.scala 31:58]
  wire [63:0] _mem_result_T_18 = {32'h0,io_cache_io_rdata_rep_bits_rdata[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _mem_result_T_19 = addr_temp[2] ? _mem_result_T_15 : _mem_result_T_18; // @[MEM.scala 154:24]
  wire [7:0] _mem_result_T_20 = _T_15 ? io_cache_io_rdata_rep_bits_rdata[63:56] : 8'h0; // @[Mux.scala 101:16]
  wire [7:0] _mem_result_T_21 = _T_13 ? io_cache_io_rdata_rep_bits_rdata[55:48] : _mem_result_T_20; // @[Mux.scala 101:16]
  wire [7:0] _mem_result_T_22 = _T_11 ? io_cache_io_rdata_rep_bits_rdata[47:40] : _mem_result_T_21; // @[Mux.scala 101:16]
  wire [7:0] _mem_result_T_23 = _T_9 ? io_cache_io_rdata_rep_bits_rdata[39:32] : _mem_result_T_22; // @[Mux.scala 101:16]
  wire [7:0] _mem_result_T_24 = _T_7 ? io_cache_io_rdata_rep_bits_rdata[31:24] : _mem_result_T_23; // @[Mux.scala 101:16]
  wire [7:0] _mem_result_T_25 = _T_5 ? io_cache_io_rdata_rep_bits_rdata[23:16] : _mem_result_T_24; // @[Mux.scala 101:16]
  wire [7:0] _mem_result_T_26 = _T_3 ? io_cache_io_rdata_rep_bits_rdata[15:8] : _mem_result_T_25; // @[Mux.scala 101:16]
  wire [7:0] _mem_result_T_27 = _T_1 ? io_cache_io_rdata_rep_bits_rdata[7:0] : _mem_result_T_26; // @[Mux.scala 101:16]
  wire [63:0] _mem_result_T_29 = {56'h0,_mem_result_T_27}; // @[Cat.scala 31:58]
  wire  mem_result_sign_2 = _mem_result_T_27[7]; // @[util.scala 11:19]
  wire [55:0] _mem_result_T_39 = mem_result_sign_2 ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _mem_result_T_40 = {_mem_result_T_39,_mem_result_T_27}; // @[Cat.scala 31:58]
  wire [15:0] _mem_result_T_41 = _T_116 ? io_cache_io_rdata_rep_bits_rdata[63:48] : 16'h0; // @[Mux.scala 101:16]
  wire [15:0] _mem_result_T_42 = _T_113 ? io_cache_io_rdata_rep_bits_rdata[47:32] : _mem_result_T_41; // @[Mux.scala 101:16]
  wire [15:0] _mem_result_T_43 = _T_110 ? io_cache_io_rdata_rep_bits_rdata[31:16] : _mem_result_T_42; // @[Mux.scala 101:16]
  wire [15:0] _mem_result_T_44 = _T_107 ? io_cache_io_rdata_rep_bits_rdata[15:0] : _mem_result_T_43; // @[Mux.scala 101:16]
  wire  mem_result_sign_3 = _mem_result_T_44[15]; // @[util.scala 11:19]
  wire [47:0] _mem_result_T_46 = mem_result_sign_3 ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _mem_result_T_47 = {_mem_result_T_46,_mem_result_T_44}; // @[Cat.scala 31:58]
  wire [63:0] _mem_result_T_53 = {48'h0,_mem_result_T_44}; // @[Cat.scala 31:58]
  wire [63:0] _GEN_36 = _T_72 ? _mem_result_T_53 : 64'h0; // @[MEM.scala 146:44 166:18]
  wire [63:0] _GEN_37 = _T_71 ? _mem_result_T_47 : _GEN_36; // @[MEM.scala 146:44 163:18]
  wire [63:0] _GEN_38 = _T_68 ? _mem_result_T_40 : _GEN_37; // @[MEM.scala 146:44 160:18]
  wire [63:0] _GEN_39 = _T_67 ? _mem_result_T_29 : _GEN_38; // @[MEM.scala 146:44 157:18]
  wire [63:0] _GEN_40 = _T_66 ? _mem_result_T_19 : _GEN_39; // @[MEM.scala 146:44 154:18]
  wire [63:0] _GEN_41 = _T_65 ? _mem_result_T_10 : _GEN_40; // @[MEM.scala 146:44 151:18]
  wire [63:0] mem_result = _T_62 ? io_cache_io_rdata_rep_bits_rdata : _GEN_41; // @[MEM.scala 146:44 148:18]
  wire  _io_out_bits_ctrl_rf_rfData_T = io_in_bits_ctrl_signal_fuType == 3'h4; // @[MEM.scala 176:67]
  wire  _io_cache_io_addr_req_valid_T_1 = _io_out_bits_ctrl_rf_rfData_T & io_in_valid; // @[MEM.scala 179:82]
  wire  _io_out_valid_T_6 = io_in_valid & _io_out_bits_ctrl_rf_rfData_T & (~io_cache_io_rdata_rep_valid & ~
    io_cache_io_wdata_rep); // @[MEM.scala 194:96]
  assign io_in_ready = _io_out_valid_T_6 ? 1'h0 : 1'h1; // @[MEM.scala 195:21]
  assign io_out_valid = ~io_in_valid | io_in_valid & _io_out_bits_ctrl_rf_rfData_T & (~io_cache_io_rdata_rep_valid & ~
    io_cache_io_wdata_rep) ? 1'h0 : 1'h1; // @[MEM.scala 194:22]
  assign io_out_bits_ctrl_signal_inst_valid = io_in_valid & io_in_bits_ctrl_signal_inst_valid; // @[MEM.scala 175:44]
  assign io_out_bits_ctrl_signal_rfWen = io_in_bits_ctrl_signal_rfWen; // @[MEM.scala 171:27]
  assign io_out_bits_ctrl_flow_PC = io_in_bits_ctrl_flow_PC; // @[MEM.scala 172:25]
  assign io_out_bits_ctrl_flow_inst = io_in_bits_ctrl_flow_inst; // @[MEM.scala 172:25]
  assign io_out_bits_ctrl_flow_Dnpc = io_in_bits_ctrl_flow_Dnpc; // @[MEM.scala 172:25]
  assign io_out_bits_ctrl_flow_skip = addr_temp == 64'ha0000048 | addr_temp == 64'ha00003f8 | addr_temp >= 64'ha0000000
     & addr_temp <= 64'ha1200000; // @[MEM.scala 174:97]
  assign io_out_bits_ctrl_rf_rfDest = io_in_bits_ctrl_rf_rfDest; // @[MEM.scala 173:23]
  assign io_out_bits_ctrl_rf_rfWen = io_in_valid & io_in_bits_ctrl_signal_rfWen; // @[MEM.scala 177:35]
  assign io_out_bits_ctrl_rf_rfData = io_in_bits_ctrl_signal_fuType == 3'h4 ? mem_result : io_in_bits_ctrl_rf_rfData; // @[MEM.scala 176:36]
  assign io_cache_io_addr_req_valid = _io_out_bits_ctrl_rf_rfData_T & io_in_valid & io_out_bits_ctrl_signal_inst_valid; // @[MEM.scala 179:97]
  assign io_cache_io_addr_req_bits_addr = 7'h45 == io_in_bits_ctrl_signal_aluoptype ? _addr_temp_T_1 : _GEN_16; // @[MEM.scala 54:44 56:17]
  assign io_cache_io_addr_req_bits_ce = _io_cache_io_addr_req_valid_T_1 & io_out_bits_ctrl_signal_inst_valid; // @[MEM.scala 181:99]
  assign io_cache_io_addr_req_bits_we = 7'h45 == io_in_bits_ctrl_signal_aluoptype ? 1'h0 : _GEN_17; // @[MEM.scala 54:44]
  assign io_cache_io_wdata_req_bits_wdata = _T_63 ? io_in_bits_ctrl_data_src2 : _GEN_33; // @[MEM.scala 93:44 97:18]
  assign io_cache_io_wdata_req_bits_wmask = _T_63 ? 8'hff : _GEN_32; // @[MEM.scala 93:44 96:18]
endmodule
module WB(
  input         io_in_valid,
  input         io_in_bits_ctrl_signal_inst_valid,
  input         io_in_bits_ctrl_signal_rfWen,
  input  [63:0] io_in_bits_ctrl_flow_PC,
  input  [31:0] io_in_bits_ctrl_flow_inst,
  input  [63:0] io_in_bits_ctrl_flow_Dnpc,
  input         io_in_bits_ctrl_flow_skip,
  input  [4:0]  io_in_bits_ctrl_rf_rfDest,
  input  [63:0] io_in_bits_ctrl_rf_rfData,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_ctrl_signal_inst_valid,
  output [63:0] io_out_bits_ctrl_flow_PC,
  output [31:0] io_out_bits_ctrl_flow_inst,
  output [63:0] io_out_bits_ctrl_flow_Dnpc,
  output        io_out_bits_ctrl_flow_skip,
  output [4:0]  io_out_bits_ctrl_rf_rfDest,
  output        io_out_bits_ctrl_rf_rfWen,
  output [63:0] io_out_bits_ctrl_rf_rfData
);
  assign io_out_valid = io_in_valid; // @[WB.scala 18:22]
  assign io_out_bits_ctrl_signal_inst_valid = io_in_valid & io_in_bits_ctrl_signal_inst_valid; // @[WB.scala 15:44]
  assign io_out_bits_ctrl_flow_PC = io_in_bits_ctrl_flow_PC; // @[WB.scala 13:15]
  assign io_out_bits_ctrl_flow_inst = io_in_bits_ctrl_flow_inst; // @[WB.scala 13:15]
  assign io_out_bits_ctrl_flow_Dnpc = io_in_bits_ctrl_flow_Dnpc; // @[WB.scala 13:15]
  assign io_out_bits_ctrl_flow_skip = io_in_bits_ctrl_flow_skip; // @[WB.scala 13:15]
  assign io_out_bits_ctrl_rf_rfDest = io_in_bits_ctrl_rf_rfDest; // @[WB.scala 13:15]
  assign io_out_bits_ctrl_rf_rfWen = io_in_valid & io_in_bits_ctrl_signal_rfWen; // @[WB.scala 16:35]
  assign io_out_bits_ctrl_rf_rfData = io_in_bits_ctrl_rf_rfData; // @[WB.scala 13:15]
endmodule
module Bypass(
  input  [4:0]  io_EX_rf_rfDest,
  input         io_EX_rf_rfWen,
  input  [63:0] io_EX_rf_rfData,
  input  [4:0]  io_MEM_rf_rfDest,
  input         io_MEM_rf_rfWen,
  input  [63:0] io_MEM_rf_rfData,
  input  [4:0]  io_WB_rf_rfDest,
  input         io_WB_rf_rfWen,
  input  [63:0] io_WB_rf_rfData,
  input  [63:0] io_Reg1,
  input  [4:0]  io_reg_index1,
  input  [63:0] io_Reg2,
  input  [4:0]  io_reg_index2,
  output [63:0] io_Bypass_REG1,
  output [63:0] io_Bypass_REG2
);
  wire  _reg1_temp_T_3 = io_EX_rf_rfDest != 5'h0; // @[Bypass.scala 26:92]
  wire  _reg1_temp_T_4 = io_EX_rf_rfWen & io_EX_rf_rfDest == io_reg_index1 & io_EX_rf_rfDest != 5'h0; // @[Bypass.scala 26:73]
  wire  _reg1_temp_T_8 = io_MEM_rf_rfDest != 5'h0; // @[Bypass.scala 27:95]
  wire  _reg1_temp_T_9 = io_MEM_rf_rfWen & io_MEM_rf_rfDest == io_reg_index1 & io_MEM_rf_rfDest != 5'h0; // @[Bypass.scala 27:75]
  wire  _reg1_temp_T_13 = io_WB_rf_rfDest != 5'h0; // @[Bypass.scala 28:92]
  wire  _reg1_temp_T_14 = io_WB_rf_rfWen & io_WB_rf_rfDest == io_reg_index1 & io_WB_rf_rfDest != 5'h0; // @[Bypass.scala 28:73]
  wire [63:0] _reg1_temp_T_15 = _reg1_temp_T_14 ? io_WB_rf_rfData : io_Reg1; // @[Mux.scala 47:70]
  wire [63:0] _reg1_temp_T_16 = _reg1_temp_T_9 ? io_MEM_rf_rfData : _reg1_temp_T_15; // @[Mux.scala 47:70]
  wire  _reg2_temp_T_4 = io_EX_rf_rfWen & io_EX_rf_rfDest == io_reg_index2 & _reg1_temp_T_3; // @[Bypass.scala 34:73]
  wire  _reg2_temp_T_9 = io_MEM_rf_rfWen & io_MEM_rf_rfDest == io_reg_index2 & _reg1_temp_T_8; // @[Bypass.scala 35:75]
  wire  _reg2_temp_T_14 = io_WB_rf_rfWen & io_WB_rf_rfDest == io_reg_index2 & _reg1_temp_T_13; // @[Bypass.scala 36:73]
  wire [63:0] _reg2_temp_T_15 = _reg2_temp_T_14 ? io_WB_rf_rfData : io_Reg2; // @[Mux.scala 47:70]
  wire [63:0] _reg2_temp_T_16 = _reg2_temp_T_9 ? io_MEM_rf_rfData : _reg2_temp_T_15; // @[Mux.scala 47:70]
  assign io_Bypass_REG1 = _reg1_temp_T_4 ? io_EX_rf_rfData : _reg1_temp_T_16; // @[Mux.scala 47:70]
  assign io_Bypass_REG2 = _reg2_temp_T_4 ? io_EX_rf_rfData : _reg2_temp_T_16; // @[Mux.scala 47:70]
endmodule
module MEM_Bypass(
  input  [4:0]  io_MEM_rf_rfDest,
  input         io_MEM_rf_rfWen,
  input  [63:0] io_MEM_rf_rfData,
  input  [63:0] io_Reg1,
  input  [4:0]  io_reg_index1,
  input  [63:0] io_Reg2,
  input  [4:0]  io_reg_index2,
  output [63:0] io_Bypass_REG1,
  output [63:0] io_Bypass_REG2
);
  wire  _reg1_temp_T_3 = io_MEM_rf_rfDest != 5'h0; // @[Bypass.scala 66:95]
  wire  _reg1_temp_T_4 = io_MEM_rf_rfWen & io_MEM_rf_rfDest == io_reg_index1 & io_MEM_rf_rfDest != 5'h0; // @[Bypass.scala 66:75]
  wire  _reg2_temp_T_4 = io_MEM_rf_rfWen & io_MEM_rf_rfDest == io_reg_index2 & _reg1_temp_T_3; // @[Bypass.scala 72:75]
  assign io_Bypass_REG1 = _reg1_temp_T_4 ? io_MEM_rf_rfData : io_Reg1; // @[Mux.scala 47:70]
  assign io_Bypass_REG2 = _reg2_temp_T_4 ? io_MEM_rf_rfData : io_Reg2; // @[Mux.scala 47:70]
endmodule
module Cache_Data(
  input          clock,
  input          io_in_valid,
  input  [63:0]  io_in_addr,
  input  [63:0]  io_write_bus_addr,
  input          io_write_bus_valid,
  input  [1:0]   io_write_bus_waymask,
  input  [511:0] io_write_bus_wdata,
  output         io_out_valid,
  output [52:0]  io_out_bits_meat_tag_0,
  output [52:0]  io_out_bits_meat_tag_1,
  output         io_out_bits_meat_valid_0,
  output         io_out_bits_meat_valid_1,
  output [511:0] io_out_bits_data_data_0,
  output [511:0] io_out_bits_data_data_1,
  output [52:0]  io_out_bits_ctrl_data_tag,
  output [4:0]   io_out_bits_ctrl_data_index,
  output [5:0]   io_out_bits_ctrl_data_offset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [511:0] _RAND_0;
  reg [511:0] _RAND_3;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  reg [511:0] data_0 [0:31]; // @[Cache.scala 119:25]
  wire  data_0_data_w_en; // @[Cache.scala 119:25]
  wire [4:0] data_0_data_w_addr; // @[Cache.scala 119:25]
  wire [511:0] data_0_data_w_data; // @[Cache.scala 119:25]
  wire [511:0] data_0_MPORT_data; // @[Cache.scala 119:25]
  wire [4:0] data_0_MPORT_addr; // @[Cache.scala 119:25]
  wire  data_0_MPORT_mask; // @[Cache.scala 119:25]
  wire  data_0_MPORT_en; // @[Cache.scala 119:25]
  reg  data_0_data_w_en_pipe_0;
  reg [4:0] data_0_data_w_addr_pipe_0;
  reg [511:0] data_1 [0:31]; // @[Cache.scala 119:25]
  wire  data_1_data_w_en; // @[Cache.scala 119:25]
  wire [4:0] data_1_data_w_addr; // @[Cache.scala 119:25]
  wire [511:0] data_1_data_w_data; // @[Cache.scala 119:25]
  wire [511:0] data_1_MPORT_data; // @[Cache.scala 119:25]
  wire [4:0] data_1_MPORT_addr; // @[Cache.scala 119:25]
  wire  data_1_MPORT_mask; // @[Cache.scala 119:25]
  wire  data_1_MPORT_en; // @[Cache.scala 119:25]
  reg  data_1_data_w_en_pipe_0;
  reg [4:0] data_1_data_w_addr_pipe_0;
  reg [52:0] TAG_0 [0:31]; // @[Cache.scala 121:24]
  wire  TAG_0_tag_w_en; // @[Cache.scala 121:24]
  wire [4:0] TAG_0_tag_w_addr; // @[Cache.scala 121:24]
  wire [52:0] TAG_0_tag_w_data; // @[Cache.scala 121:24]
  wire [52:0] TAG_0_MPORT_1_data; // @[Cache.scala 121:24]
  wire [4:0] TAG_0_MPORT_1_addr; // @[Cache.scala 121:24]
  wire  TAG_0_MPORT_1_mask; // @[Cache.scala 121:24]
  wire  TAG_0_MPORT_1_en; // @[Cache.scala 121:24]
  reg  TAG_0_tag_w_en_pipe_0;
  reg [4:0] TAG_0_tag_w_addr_pipe_0;
  reg [52:0] TAG_1 [0:31]; // @[Cache.scala 121:24]
  wire  TAG_1_tag_w_en; // @[Cache.scala 121:24]
  wire [4:0] TAG_1_tag_w_addr; // @[Cache.scala 121:24]
  wire [52:0] TAG_1_tag_w_data; // @[Cache.scala 121:24]
  wire [52:0] TAG_1_MPORT_1_data; // @[Cache.scala 121:24]
  wire [4:0] TAG_1_MPORT_1_addr; // @[Cache.scala 121:24]
  wire  TAG_1_MPORT_1_mask; // @[Cache.scala 121:24]
  wire  TAG_1_MPORT_1_en; // @[Cache.scala 121:24]
  reg  TAG_1_tag_w_en_pipe_0;
  reg [4:0] TAG_1_tag_w_addr_pipe_0;
  reg  data_valid_0 [0:31]; // @[Cache.scala 122:31]
  wire  data_valid_0_valid_w_en; // @[Cache.scala 122:31]
  wire [4:0] data_valid_0_valid_w_addr; // @[Cache.scala 122:31]
  wire  data_valid_0_valid_w_data; // @[Cache.scala 122:31]
  wire  data_valid_0_MPORT_2_data; // @[Cache.scala 122:31]
  wire [4:0] data_valid_0_MPORT_2_addr; // @[Cache.scala 122:31]
  wire  data_valid_0_MPORT_2_mask; // @[Cache.scala 122:31]
  wire  data_valid_0_MPORT_2_en; // @[Cache.scala 122:31]
  reg  data_valid_0_valid_w_en_pipe_0;
  reg [4:0] data_valid_0_valid_w_addr_pipe_0;
  reg  data_valid_1 [0:31]; // @[Cache.scala 122:31]
  wire  data_valid_1_valid_w_en; // @[Cache.scala 122:31]
  wire [4:0] data_valid_1_valid_w_addr; // @[Cache.scala 122:31]
  wire  data_valid_1_valid_w_data; // @[Cache.scala 122:31]
  wire  data_valid_1_MPORT_2_data; // @[Cache.scala 122:31]
  wire [4:0] data_valid_1_MPORT_2_addr; // @[Cache.scala 122:31]
  wire  data_valid_1_MPORT_2_mask; // @[Cache.scala 122:31]
  wire  data_valid_1_MPORT_2_en; // @[Cache.scala 122:31]
  reg  data_valid_1_valid_w_en_pipe_0;
  reg [4:0] data_valid_1_valid_w_addr_pipe_0;
  assign data_0_data_w_en = data_0_data_w_en_pipe_0;
  assign data_0_data_w_addr = data_0_data_w_addr_pipe_0;
  assign data_0_data_w_data = data_0[data_0_data_w_addr]; // @[Cache.scala 119:25]
  assign data_0_MPORT_data = io_write_bus_wdata;
  assign data_0_MPORT_addr = io_write_bus_addr[10:6];
  assign data_0_MPORT_mask = io_write_bus_waymask[0];
  assign data_0_MPORT_en = io_write_bus_valid;
  assign data_1_data_w_en = data_1_data_w_en_pipe_0;
  assign data_1_data_w_addr = data_1_data_w_addr_pipe_0;
  assign data_1_data_w_data = data_1[data_1_data_w_addr]; // @[Cache.scala 119:25]
  assign data_1_MPORT_data = io_write_bus_wdata;
  assign data_1_MPORT_addr = io_write_bus_addr[10:6];
  assign data_1_MPORT_mask = io_write_bus_waymask[1];
  assign data_1_MPORT_en = io_write_bus_valid;
  assign TAG_0_tag_w_en = TAG_0_tag_w_en_pipe_0;
  assign TAG_0_tag_w_addr = TAG_0_tag_w_addr_pipe_0;
  assign TAG_0_tag_w_data = TAG_0[TAG_0_tag_w_addr]; // @[Cache.scala 121:24]
  assign TAG_0_MPORT_1_data = io_write_bus_addr[63:11];
  assign TAG_0_MPORT_1_addr = io_write_bus_addr[10:6];
  assign TAG_0_MPORT_1_mask = io_write_bus_waymask[0];
  assign TAG_0_MPORT_1_en = io_write_bus_valid;
  assign TAG_1_tag_w_en = TAG_1_tag_w_en_pipe_0;
  assign TAG_1_tag_w_addr = TAG_1_tag_w_addr_pipe_0;
  assign TAG_1_tag_w_data = TAG_1[TAG_1_tag_w_addr]; // @[Cache.scala 121:24]
  assign TAG_1_MPORT_1_data = io_write_bus_addr[63:11];
  assign TAG_1_MPORT_1_addr = io_write_bus_addr[10:6];
  assign TAG_1_MPORT_1_mask = io_write_bus_waymask[1];
  assign TAG_1_MPORT_1_en = io_write_bus_valid;
  assign data_valid_0_valid_w_en = data_valid_0_valid_w_en_pipe_0;
  assign data_valid_0_valid_w_addr = data_valid_0_valid_w_addr_pipe_0;
  assign data_valid_0_valid_w_data = data_valid_0[data_valid_0_valid_w_addr]; // @[Cache.scala 122:31]
  assign data_valid_0_MPORT_2_data = 1'h1;
  assign data_valid_0_MPORT_2_addr = io_write_bus_addr[10:6];
  assign data_valid_0_MPORT_2_mask = io_write_bus_waymask[0];
  assign data_valid_0_MPORT_2_en = io_write_bus_valid;
  assign data_valid_1_valid_w_en = data_valid_1_valid_w_en_pipe_0;
  assign data_valid_1_valid_w_addr = data_valid_1_valid_w_addr_pipe_0;
  assign data_valid_1_valid_w_data = data_valid_1[data_valid_1_valid_w_addr]; // @[Cache.scala 122:31]
  assign data_valid_1_MPORT_2_data = 1'h1;
  assign data_valid_1_MPORT_2_addr = io_write_bus_addr[10:6];
  assign data_valid_1_MPORT_2_mask = io_write_bus_waymask[1];
  assign data_valid_1_MPORT_2_en = io_write_bus_valid;
  assign io_out_valid = io_in_valid; // @[Cache.scala 138:22]
  assign io_out_bits_meat_tag_0 = TAG_0_tag_w_data; // @[Cache.scala 136:24]
  assign io_out_bits_meat_tag_1 = TAG_1_tag_w_data; // @[Cache.scala 136:24]
  assign io_out_bits_meat_valid_0 = data_valid_0_valid_w_data; // @[Cache.scala 133:26]
  assign io_out_bits_meat_valid_1 = data_valid_1_valid_w_data; // @[Cache.scala 133:26]
  assign io_out_bits_data_data_0 = data_0_data_w_data; // @[Cache.scala 134:25]
  assign io_out_bits_data_data_1 = data_1_data_w_data; // @[Cache.scala 134:25]
  assign io_out_bits_ctrl_data_tag = io_in_addr[63:11]; // @[Cache.scala 114:23]
  assign io_out_bits_ctrl_data_index = io_in_addr[10:6]; // @[Cache.scala 115:25]
  assign io_out_bits_ctrl_data_offset = io_in_addr[5:0]; // @[Cache.scala 116:26]
  always @(posedge clock) begin
    if (data_0_MPORT_en & data_0_MPORT_mask) begin
      data_0[data_0_MPORT_addr] <= data_0_MPORT_data; // @[Cache.scala 119:25]
    end
    data_0_data_w_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      data_0_data_w_addr_pipe_0 <= io_in_addr[10:6];
    end
    if (data_1_MPORT_en & data_1_MPORT_mask) begin
      data_1[data_1_MPORT_addr] <= data_1_MPORT_data; // @[Cache.scala 119:25]
    end
    data_1_data_w_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      data_1_data_w_addr_pipe_0 <= io_in_addr[10:6];
    end
    if (TAG_0_MPORT_1_en & TAG_0_MPORT_1_mask) begin
      TAG_0[TAG_0_MPORT_1_addr] <= TAG_0_MPORT_1_data; // @[Cache.scala 121:24]
    end
    TAG_0_tag_w_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      TAG_0_tag_w_addr_pipe_0 <= io_in_addr[10:6];
    end
    if (TAG_1_MPORT_1_en & TAG_1_MPORT_1_mask) begin
      TAG_1[TAG_1_MPORT_1_addr] <= TAG_1_MPORT_1_data; // @[Cache.scala 121:24]
    end
    TAG_1_tag_w_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      TAG_1_tag_w_addr_pipe_0 <= io_in_addr[10:6];
    end
    if (data_valid_0_MPORT_2_en & data_valid_0_MPORT_2_mask) begin
      data_valid_0[data_valid_0_MPORT_2_addr] <= data_valid_0_MPORT_2_data; // @[Cache.scala 122:31]
    end
    data_valid_0_valid_w_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      data_valid_0_valid_w_addr_pipe_0 <= io_in_addr[10:6];
    end
    if (data_valid_1_MPORT_2_en & data_valid_1_MPORT_2_mask) begin
      data_valid_1[data_valid_1_MPORT_2_addr] <= data_valid_1_MPORT_2_data; // @[Cache.scala 122:31]
    end
    data_valid_1_valid_w_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      data_valid_1_valid_w_addr_pipe_0 <= io_in_addr[10:6];
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {16{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    data_0[initvar] = _RAND_0[511:0];
  _RAND_3 = {16{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    data_1[initvar] = _RAND_3[511:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    TAG_0[initvar] = _RAND_6[52:0];
  _RAND_9 = {2{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    TAG_1[initvar] = _RAND_9[52:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    data_valid_0[initvar] = _RAND_12[0:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    data_valid_1[initvar] = _RAND_15[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  data_0_data_w_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_data_w_addr_pipe_0 = _RAND_2[4:0];
  _RAND_4 = {1{`RANDOM}};
  data_1_data_w_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  data_1_data_w_addr_pipe_0 = _RAND_5[4:0];
  _RAND_7 = {1{`RANDOM}};
  TAG_0_tag_w_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  TAG_0_tag_w_addr_pipe_0 = _RAND_8[4:0];
  _RAND_10 = {1{`RANDOM}};
  TAG_1_tag_w_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  TAG_1_tag_w_addr_pipe_0 = _RAND_11[4:0];
  _RAND_13 = {1{`RANDOM}};
  data_valid_0_valid_w_en_pipe_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  data_valid_0_valid_w_addr_pipe_0 = _RAND_14[4:0];
  _RAND_16 = {1{`RANDOM}};
  data_valid_1_valid_w_en_pipe_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  data_valid_1_valid_w_addr_pipe_0 = _RAND_17[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scanf_data(
  input          io_in_valid,
  input  [52:0]  io_in_bits_meat_tag_0,
  input  [52:0]  io_in_bits_meat_tag_1,
  input          io_in_bits_meat_valid_0,
  input          io_in_bits_meat_valid_1,
  input  [511:0] io_in_bits_data_data_0,
  input  [511:0] io_in_bits_data_data_1,
  input  [52:0]  io_in_bits_ctrl_data_tag,
  input  [4:0]   io_in_bits_ctrl_data_index,
  output         io_out_bits_hit,
  output [511:0] io_out_bits_data,
  output [4:0]   io_out_bits_meta_ctrl_data_index,
  output         io_out_bits_hit_way_0,
  output         io_out_bits_hit_way_1,
  output [52:0]  io_out_bits_tag_0,
  output [52:0]  io_out_bits_tag_1
);
  wire  _hit_way_0_T = io_in_bits_meat_valid_0 & io_in_valid; // @[Cache.scala 74:98]
  wire  hit_way_0_result = _hit_way_0_T & io_in_bits_ctrl_data_tag == io_in_bits_meat_tag_0; // @[Cache.scala 68:20]
  wire  _hit_way_1_T = io_in_bits_meat_valid_1 & io_in_valid; // @[Cache.scala 74:98]
  wire  hit_way_1_result = _hit_way_1_T & io_in_bits_ctrl_data_tag == io_in_bits_meat_tag_1; // @[Cache.scala 68:20]
  wire [511:0] _GEN_3 = hit_way_0_result ? io_in_bits_data_data_0 : 512'h0; // @[Cache.scala 80:29 82:17]
  assign io_out_bits_hit = hit_way_1_result | hit_way_0_result; // @[Cache.scala 80:29 81:16]
  assign io_out_bits_data = hit_way_1_result ? io_in_bits_data_data_1 : _GEN_3; // @[Cache.scala 80:29 82:17]
  assign io_out_bits_meta_ctrl_data_index = io_in_bits_ctrl_data_index; // @[Cache.scala 90:30]
  assign io_out_bits_hit_way_0 = _hit_way_0_T & io_in_bits_ctrl_data_tag == io_in_bits_meat_tag_0; // @[Cache.scala 68:20]
  assign io_out_bits_hit_way_1 = _hit_way_1_T & io_in_bits_ctrl_data_tag == io_in_bits_meat_tag_1; // @[Cache.scala 68:20]
  assign io_out_bits_tag_0 = io_in_bits_meat_tag_0; // @[Cache.scala 96:19]
  assign io_out_bits_tag_1 = io_in_bits_meat_tag_1; // @[Cache.scala 96:19]
endmodule
module Cache(
  input         clock,
  input         reset,
  input         io_in_addr_req_valid,
  input  [63:0] io_in_addr_req_bits_addr,
  input         io_in_rdata_rep_ready,
  output        io_in_rdata_rep_valid,
  output [63:0] io_in_rdata_rep_bits_rdata,
  input         io_flush,
  output        io_out_addr_req_valid,
  output [63:0] io_out_addr_req_bits_addr,
  output        io_out_addr_req_bits_ce,
  input         io_out_rdata_rep_valid,
  input  [63:0] io_out_rdata_rep_bits_rdata
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [511:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  Cache_data_clock; // @[Cache.scala 159:26]
  wire  Cache_data_io_in_valid; // @[Cache.scala 159:26]
  wire [63:0] Cache_data_io_in_addr; // @[Cache.scala 159:26]
  wire [63:0] Cache_data_io_write_bus_addr; // @[Cache.scala 159:26]
  wire  Cache_data_io_write_bus_valid; // @[Cache.scala 159:26]
  wire [1:0] Cache_data_io_write_bus_waymask; // @[Cache.scala 159:26]
  wire [511:0] Cache_data_io_write_bus_wdata; // @[Cache.scala 159:26]
  wire  Cache_data_io_out_valid; // @[Cache.scala 159:26]
  wire [52:0] Cache_data_io_out_bits_meat_tag_0; // @[Cache.scala 159:26]
  wire [52:0] Cache_data_io_out_bits_meat_tag_1; // @[Cache.scala 159:26]
  wire  Cache_data_io_out_bits_meat_valid_0; // @[Cache.scala 159:26]
  wire  Cache_data_io_out_bits_meat_valid_1; // @[Cache.scala 159:26]
  wire [511:0] Cache_data_io_out_bits_data_data_0; // @[Cache.scala 159:26]
  wire [511:0] Cache_data_io_out_bits_data_data_1; // @[Cache.scala 159:26]
  wire [52:0] Cache_data_io_out_bits_ctrl_data_tag; // @[Cache.scala 159:26]
  wire [4:0] Cache_data_io_out_bits_ctrl_data_index; // @[Cache.scala 159:26]
  wire [5:0] Cache_data_io_out_bits_ctrl_data_offset; // @[Cache.scala 159:26]
  wire  Scanf_io_in_valid; // @[Cache.scala 160:21]
  wire [52:0] Scanf_io_in_bits_meat_tag_0; // @[Cache.scala 160:21]
  wire [52:0] Scanf_io_in_bits_meat_tag_1; // @[Cache.scala 160:21]
  wire  Scanf_io_in_bits_meat_valid_0; // @[Cache.scala 160:21]
  wire  Scanf_io_in_bits_meat_valid_1; // @[Cache.scala 160:21]
  wire [511:0] Scanf_io_in_bits_data_data_0; // @[Cache.scala 160:21]
  wire [511:0] Scanf_io_in_bits_data_data_1; // @[Cache.scala 160:21]
  wire [52:0] Scanf_io_in_bits_ctrl_data_tag; // @[Cache.scala 160:21]
  wire [4:0] Scanf_io_in_bits_ctrl_data_index; // @[Cache.scala 160:21]
  wire  Scanf_io_out_bits_hit; // @[Cache.scala 160:21]
  wire [511:0] Scanf_io_out_bits_data; // @[Cache.scala 160:21]
  wire [4:0] Scanf_io_out_bits_meta_ctrl_data_index; // @[Cache.scala 160:21]
  wire  Scanf_io_out_bits_hit_way_0; // @[Cache.scala 160:21]
  wire  Scanf_io_out_bits_hit_way_1; // @[Cache.scala 160:21]
  wire [52:0] Scanf_io_out_bits_tag_0; // @[Cache.scala 160:21]
  wire [52:0] Scanf_io_out_bits_tag_1; // @[Cache.scala 160:21]
  reg  lru [0:31]; // @[Cache.scala 173:24]
  wire  lru_lru_w_MPORT_en; // @[Cache.scala 173:24]
  wire [4:0] lru_lru_w_MPORT_addr; // @[Cache.scala 173:24]
  wire  lru_lru_w_MPORT_data; // @[Cache.scala 173:24]
  wire  lru_MPORT_data; // @[Cache.scala 173:24]
  wire [4:0] lru_MPORT_addr; // @[Cache.scala 173:24]
  wire  lru_MPORT_mask; // @[Cache.scala 173:24]
  wire  lru_MPORT_en; // @[Cache.scala 173:24]
  wire  lru_MPORT_1_data; // @[Cache.scala 173:24]
  wire [4:0] lru_MPORT_1_addr; // @[Cache.scala 173:24]
  wire  lru_MPORT_1_mask; // @[Cache.scala 173:24]
  wire  lru_MPORT_1_en; // @[Cache.scala 173:24]
  wire  lru_MPORT_2_data; // @[Cache.scala 173:24]
  wire [4:0] lru_MPORT_2_addr; // @[Cache.scala 173:24]
  wire  lru_MPORT_2_mask; // @[Cache.scala 173:24]
  wire  lru_MPORT_2_en; // @[Cache.scala 173:24]
  wire  lru_MPORT_3_data; // @[Cache.scala 173:24]
  wire [4:0] lru_MPORT_3_addr; // @[Cache.scala 173:24]
  wire  lru_MPORT_3_mask; // @[Cache.scala 173:24]
  wire  lru_MPORT_3_en; // @[Cache.scala 173:24]
  reg  lru_lru_w_MPORT_en_pipe_0;
  reg [4:0] lru_lru_w_MPORT_addr_pipe_0;
  reg [1:0] state; // @[Cache.scala 163:22]
  reg [511:0] data_line_reg; // @[Cache.scala 165:30]
  reg [63:0] mem_addr_reg; // @[Cache.scala 166:29]
  reg  lru_r; // @[Cache.scala 168:23]
  reg [3:0] count; // @[Cache.scala 176:22]
  wire  s = count == 4'h8; // @[Cache.scala 177:17]
  wire  _T = 2'h0 == state; // @[Cache.scala 196:16]
  wire  _T_1 = 2'h1 == state; // @[Cache.scala 196:16]
  wire [63:0] _mem_addr_reg_T_2 = {io_in_addr_req_bits_addr[63:6],6'h0}; // @[Cat.scala 31:58]
  wire  hit_way_0 = Scanf_io_out_bits_hit_way_0; // @[Cache.scala 192:21 357:11]
  wire  hit_way_1 = Scanf_io_out_bits_hit_way_1; // @[Cache.scala 192:21 357:11]
  wire  lru_w = lru_lru_w_MPORT_data;
  wire  _GEN_17 = ~Scanf_io_out_bits_hit ? 1'h0 : hit_way_0; // @[Cache.scala 173:24 201:26]
  wire  _GEN_21 = ~Scanf_io_out_bits_hit ? 1'h0 : hit_way_1; // @[Cache.scala 173:24 201:26]
  wire  _T_5 = 2'h2 == state; // @[Cache.scala 196:16]
  wire [3:0] _count_T_1 = count + 4'h1; // @[Cache.scala 229:24]
  wire [63:0] _mem_addr_reg_T_4 = mem_addr_reg + 64'h8; // @[Cache.scala 230:38]
  wire [3:0] _GEN_24 = ~io_in_rdata_rep_ready & s | ~io_out_rdata_rep_valid ? count : _count_T_1; // @[Cache.scala 226:83 227:15 229:15]
  wire [63:0] _GEN_25 = ~io_in_rdata_rep_ready & s | ~io_out_rdata_rep_valid ? mem_addr_reg : _mem_addr_reg_T_4; // @[Cache.scala 166:29 226:83 230:22]
  wire [511:0] _data_line_reg_T_1 = {io_out_rdata_rep_bits_rdata,data_line_reg[511:64]}; // @[Cat.scala 31:58]
  wire [511:0] _GEN_26 = ~s & io_out_rdata_rep_valid ? _data_line_reg_T_1 : data_line_reg; // @[Cache.scala 236:51 237:23 165:30]
  wire  _GEN_34 = lru_r ? 1'h0 : 1'h1; // @[Cache.scala 173:24 240:29]
  wire  _GEN_38 = io_in_rdata_rep_ready & s & lru_r; // @[Cache.scala 173:24 239:51]
  wire  _GEN_43 = io_in_rdata_rep_ready & s & _GEN_34; // @[Cache.scala 173:24 239:51]
  wire [3:0] _GEN_45 = io_in_rdata_rep_ready & s ? 4'h0 : _GEN_24; // @[Cache.scala 239:51 245:14]
  wire  _GEN_62 = 2'h1 == state & _GEN_17; // @[Cache.scala 196:16 173:24]
  wire  _GEN_66 = 2'h1 == state & _GEN_21; // @[Cache.scala 196:16 173:24]
  wire  _GEN_73 = 2'h1 == state ? 1'h0 : 2'h2 == state & _GEN_38; // @[Cache.scala 196:16 173:24]
  wire  _GEN_78 = 2'h1 == state ? 1'h0 : 2'h2 == state & _GEN_43; // @[Cache.scala 196:16 173:24]
  wire [63:0] _GEN_102 = 3'h7 == io_in_addr_req_bits_addr[5:3] ? Scanf_io_out_bits_data[511:448] : 64'h0; // @[Cache.scala 266:115 296:16]
  wire [63:0] _GEN_103 = 3'h7 == io_in_addr_req_bits_addr[5:3] ? data_line_reg[511:448] : 64'h0; // @[Cache.scala 266:115 297:16]
  wire [63:0] _GEN_104 = 3'h6 == io_in_addr_req_bits_addr[5:3] ? Scanf_io_out_bits_data[447:384] : _GEN_102; // @[Cache.scala 266:115 292:16]
  wire [63:0] _GEN_105 = 3'h6 == io_in_addr_req_bits_addr[5:3] ? data_line_reg[447:384] : _GEN_103; // @[Cache.scala 266:115 293:16]
  wire [63:0] _GEN_106 = 3'h5 == io_in_addr_req_bits_addr[5:3] ? Scanf_io_out_bits_data[383:320] : _GEN_104; // @[Cache.scala 266:115 288:16]
  wire [63:0] _GEN_107 = 3'h5 == io_in_addr_req_bits_addr[5:3] ? data_line_reg[383:320] : _GEN_105; // @[Cache.scala 266:115 289:16]
  wire [63:0] _GEN_108 = 3'h4 == io_in_addr_req_bits_addr[5:3] ? Scanf_io_out_bits_data[319:256] : _GEN_106; // @[Cache.scala 266:115 284:16]
  wire [63:0] _GEN_109 = 3'h4 == io_in_addr_req_bits_addr[5:3] ? data_line_reg[319:256] : _GEN_107; // @[Cache.scala 266:115 285:16]
  wire [63:0] _GEN_110 = 3'h3 == io_in_addr_req_bits_addr[5:3] ? Scanf_io_out_bits_data[255:192] : _GEN_108; // @[Cache.scala 266:115 280:16]
  wire [63:0] _GEN_111 = 3'h3 == io_in_addr_req_bits_addr[5:3] ? data_line_reg[255:192] : _GEN_109; // @[Cache.scala 266:115 281:16]
  wire [63:0] _GEN_112 = 3'h2 == io_in_addr_req_bits_addr[5:3] ? Scanf_io_out_bits_data[191:128] : _GEN_110; // @[Cache.scala 266:115 276:16]
  wire [63:0] _GEN_113 = 3'h2 == io_in_addr_req_bits_addr[5:3] ? data_line_reg[191:128] : _GEN_111; // @[Cache.scala 266:115 277:16]
  wire [63:0] _GEN_114 = 3'h1 == io_in_addr_req_bits_addr[5:3] ? Scanf_io_out_bits_data[127:64] : _GEN_112; // @[Cache.scala 266:115 272:16]
  wire [63:0] _GEN_115 = 3'h1 == io_in_addr_req_bits_addr[5:3] ? data_line_reg[127:64] : _GEN_113; // @[Cache.scala 266:115 273:16]
  wire [63:0] hit_data = 3'h0 == io_in_addr_req_bits_addr[5:3] ? Scanf_io_out_bits_data[63:0] : _GEN_114; // @[Cache.scala 266:115 268:16]
  wire [63:0] mem_data = 3'h0 == io_in_addr_req_bits_addr[5:3] ? data_line_reg[63:0] : _GEN_115; // @[Cache.scala 266:115 269:16]
  wire [1:0] _GEN_119 = Scanf_io_out_bits_hit ? 2'h0 : 2'h2; // @[Cache.scala 310:26 311:17 321:19]
  wire [1:0] _GEN_120 = s & io_in_rdata_rep_ready ? 2'h0 : state; // @[Cache.scala 327:52 328:17 163:22]
  wire [1:0] _GEN_121 = _T_5 ? _GEN_120 : state; // @[Cache.scala 301:16 163:22]
  wire  _io_in_rdata_rep_bits_rdata_T_1 = state == 2'h1 & Scanf_io_out_bits_hit; // @[Cache.scala 345:54]
  reg  Scanf_io_in_valid_REG; // @[Cache.scala 352:31]
  wire  _io_out_addr_req_valid_T = state == 2'h2; // @[Cache.scala 372:40]
  wire  _io_in_rdata_rep_valid_T_4 = _io_out_addr_req_valid_T & s; // @[Cache.scala 381:75]
  Cache_Data Cache_data ( // @[Cache.scala 159:26]
    .clock(Cache_data_clock),
    .io_in_valid(Cache_data_io_in_valid),
    .io_in_addr(Cache_data_io_in_addr),
    .io_write_bus_addr(Cache_data_io_write_bus_addr),
    .io_write_bus_valid(Cache_data_io_write_bus_valid),
    .io_write_bus_waymask(Cache_data_io_write_bus_waymask),
    .io_write_bus_wdata(Cache_data_io_write_bus_wdata),
    .io_out_valid(Cache_data_io_out_valid),
    .io_out_bits_meat_tag_0(Cache_data_io_out_bits_meat_tag_0),
    .io_out_bits_meat_tag_1(Cache_data_io_out_bits_meat_tag_1),
    .io_out_bits_meat_valid_0(Cache_data_io_out_bits_meat_valid_0),
    .io_out_bits_meat_valid_1(Cache_data_io_out_bits_meat_valid_1),
    .io_out_bits_data_data_0(Cache_data_io_out_bits_data_data_0),
    .io_out_bits_data_data_1(Cache_data_io_out_bits_data_data_1),
    .io_out_bits_ctrl_data_tag(Cache_data_io_out_bits_ctrl_data_tag),
    .io_out_bits_ctrl_data_index(Cache_data_io_out_bits_ctrl_data_index),
    .io_out_bits_ctrl_data_offset(Cache_data_io_out_bits_ctrl_data_offset)
  );
  Scanf_data Scanf ( // @[Cache.scala 160:21]
    .io_in_valid(Scanf_io_in_valid),
    .io_in_bits_meat_tag_0(Scanf_io_in_bits_meat_tag_0),
    .io_in_bits_meat_tag_1(Scanf_io_in_bits_meat_tag_1),
    .io_in_bits_meat_valid_0(Scanf_io_in_bits_meat_valid_0),
    .io_in_bits_meat_valid_1(Scanf_io_in_bits_meat_valid_1),
    .io_in_bits_data_data_0(Scanf_io_in_bits_data_data_0),
    .io_in_bits_data_data_1(Scanf_io_in_bits_data_data_1),
    .io_in_bits_ctrl_data_tag(Scanf_io_in_bits_ctrl_data_tag),
    .io_in_bits_ctrl_data_index(Scanf_io_in_bits_ctrl_data_index),
    .io_out_bits_hit(Scanf_io_out_bits_hit),
    .io_out_bits_data(Scanf_io_out_bits_data),
    .io_out_bits_meta_ctrl_data_index(Scanf_io_out_bits_meta_ctrl_data_index),
    .io_out_bits_hit_way_0(Scanf_io_out_bits_hit_way_0),
    .io_out_bits_hit_way_1(Scanf_io_out_bits_hit_way_1),
    .io_out_bits_tag_0(Scanf_io_out_bits_tag_0),
    .io_out_bits_tag_1(Scanf_io_out_bits_tag_1)
  );
  assign lru_lru_w_MPORT_en = lru_lru_w_MPORT_en_pipe_0;
  assign lru_lru_w_MPORT_addr = lru_lru_w_MPORT_addr_pipe_0;
  assign lru_lru_w_MPORT_data = lru[lru_lru_w_MPORT_addr]; // @[Cache.scala 173:24]
  assign lru_MPORT_data = 1'h1;
  assign lru_MPORT_addr = Cache_data_io_out_bits_ctrl_data_index;
  assign lru_MPORT_mask = 1'h1;
  assign lru_MPORT_en = _T ? 1'h0 : _GEN_62;
  assign lru_MPORT_1_data = 1'h0;
  assign lru_MPORT_1_addr = Cache_data_io_out_bits_ctrl_data_index;
  assign lru_MPORT_1_mask = 1'h1;
  assign lru_MPORT_1_en = _T ? 1'h0 : _GEN_66;
  assign lru_MPORT_2_data = 1'h0;
  assign lru_MPORT_2_addr = Cache_data_io_out_bits_ctrl_data_index;
  assign lru_MPORT_2_mask = 1'h1;
  assign lru_MPORT_2_en = _T ? 1'h0 : _GEN_73;
  assign lru_MPORT_3_data = 1'h1;
  assign lru_MPORT_3_addr = Cache_data_io_out_bits_ctrl_data_index;
  assign lru_MPORT_3_mask = 1'h1;
  assign lru_MPORT_3_en = _T ? 1'h0 : _GEN_78;
  assign io_in_rdata_rep_valid = (_io_in_rdata_rep_bits_rdata_T_1 | _io_out_addr_req_valid_T & s) & ~io_flush; // @[Cache.scala 381:93]
  assign io_in_rdata_rep_bits_rdata = state == 2'h1 & Scanf_io_out_bits_hit ? hit_data : mem_data; // @[Cache.scala 345:36]
  assign io_out_addr_req_valid = state == 2'h2; // @[Cache.scala 372:40]
  assign io_out_addr_req_bits_addr = mem_addr_reg; // @[Cache.scala 374:31]
  assign io_out_addr_req_bits_ce = state == 2'h2; // @[Cache.scala 373:42]
  assign Cache_data_clock = clock;
  assign Cache_data_io_in_valid = io_in_addr_req_valid & state == 2'h0; // @[Cache.scala 350:54]
  assign Cache_data_io_in_addr = io_in_addr_req_bits_addr; // @[Cache.scala 351:25]
  assign Cache_data_io_write_bus_addr = _io_in_rdata_rep_valid_T_4 ? io_in_addr_req_bits_addr : 64'h0; // @[Cache.scala 418:40]
  assign Cache_data_io_write_bus_valid = count == 4'h8; // @[Cache.scala 177:17]
  assign Cache_data_io_write_bus_waymask = lru_r ? 2'h2 : 2'h1; // @[Cache.scala 420:22]
  assign Cache_data_io_write_bus_wdata = _io_in_rdata_rep_valid_T_4 ? data_line_reg : 512'h0; // @[Cache.scala 419:41]
  assign Scanf_io_in_valid = Scanf_io_in_valid_REG; // @[Cache.scala 352:21]
  assign Scanf_io_in_bits_meat_tag_0 = Cache_data_io_out_bits_meat_tag_0; // @[Cache.scala 353:25]
  assign Scanf_io_in_bits_meat_tag_1 = Cache_data_io_out_bits_meat_tag_1; // @[Cache.scala 353:25]
  assign Scanf_io_in_bits_meat_valid_0 = Cache_data_io_out_bits_meat_valid_0; // @[Cache.scala 353:25]
  assign Scanf_io_in_bits_meat_valid_1 = Cache_data_io_out_bits_meat_valid_1; // @[Cache.scala 353:25]
  assign Scanf_io_in_bits_data_data_0 = Cache_data_io_out_bits_data_data_0; // @[Cache.scala 354:25]
  assign Scanf_io_in_bits_data_data_1 = Cache_data_io_out_bits_data_data_1; // @[Cache.scala 354:25]
  assign Scanf_io_in_bits_ctrl_data_tag = Cache_data_io_out_bits_ctrl_data_tag; // @[Cache.scala 355:30]
  assign Scanf_io_in_bits_ctrl_data_index = Cache_data_io_out_bits_ctrl_data_index; // @[Cache.scala 355:30]
  always @(posedge clock) begin
    if (lru_MPORT_en & lru_MPORT_mask) begin
      lru[lru_MPORT_addr] <= lru_MPORT_data; // @[Cache.scala 173:24]
    end
    if (lru_MPORT_1_en & lru_MPORT_1_mask) begin
      lru[lru_MPORT_1_addr] <= lru_MPORT_1_data; // @[Cache.scala 173:24]
    end
    if (lru_MPORT_2_en & lru_MPORT_2_mask) begin
      lru[lru_MPORT_2_addr] <= lru_MPORT_2_data; // @[Cache.scala 173:24]
    end
    if (lru_MPORT_3_en & lru_MPORT_3_mask) begin
      lru[lru_MPORT_3_addr] <= lru_MPORT_3_data; // @[Cache.scala 173:24]
    end
    lru_lru_w_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      lru_lru_w_MPORT_addr_pipe_0 <= Cache_data_io_out_bits_ctrl_data_index;
    end
    if (reset) begin // @[Cache.scala 163:22]
      state <= 2'h0; // @[Cache.scala 163:22]
    end else if (io_flush) begin // @[Cache.scala 340:18]
      state <= 2'h0; // @[Cache.scala 341:11]
    end else if (_T) begin // @[Cache.scala 301:16]
      if (io_in_addr_req_valid) begin // @[Cache.scala 303:33]
        state <= 2'h1; // @[Cache.scala 304:15]
      end else begin
        state <= 2'h0; // @[Cache.scala 306:15]
      end
    end else if (_T_1) begin // @[Cache.scala 301:16]
      state <= _GEN_119;
    end else begin
      state <= _GEN_121;
    end
    if (reset) begin // @[Cache.scala 165:30]
      data_line_reg <= 512'h0; // @[Cache.scala 165:30]
    end else if (!(2'h0 == state)) begin // @[Cache.scala 196:16]
      if (!(2'h1 == state)) begin // @[Cache.scala 196:16]
        if (2'h2 == state) begin // @[Cache.scala 196:16]
          data_line_reg <= _GEN_26;
        end
      end
    end
    if (reset) begin // @[Cache.scala 166:29]
      mem_addr_reg <= 64'h0; // @[Cache.scala 166:29]
    end else if (!(2'h0 == state)) begin // @[Cache.scala 196:16]
      if (2'h1 == state) begin // @[Cache.scala 196:16]
        if (~Scanf_io_out_bits_hit) begin // @[Cache.scala 201:26]
          mem_addr_reg <= _mem_addr_reg_T_2; // @[Cache.scala 202:24]
        end
      end else if (2'h2 == state) begin // @[Cache.scala 196:16]
        mem_addr_reg <= _GEN_25;
      end
    end
    if (reset) begin // @[Cache.scala 168:23]
      lru_r <= 1'h0; // @[Cache.scala 168:23]
    end else if (!(2'h0 == state)) begin // @[Cache.scala 196:16]
      if (2'h1 == state) begin // @[Cache.scala 196:16]
        if (~Scanf_io_out_bits_hit) begin // @[Cache.scala 201:26]
          lru_r <= lru_w; // @[Cache.scala 203:17]
        end
      end
    end
    if (reset) begin // @[Cache.scala 176:22]
      count <= 4'h0; // @[Cache.scala 176:22]
    end else if (2'h0 == state) begin // @[Cache.scala 196:16]
      count <= 4'h0; // @[Cache.scala 198:13]
    end else if (!(2'h1 == state)) begin // @[Cache.scala 196:16]
      if (2'h2 == state) begin // @[Cache.scala 196:16]
        count <= _GEN_45;
      end
    end
    Scanf_io_in_valid_REG <= Cache_data_io_out_valid; // @[Cache.scala 352:31]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    lru[initvar] = _RAND_0[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  lru_lru_w_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  lru_lru_w_MPORT_addr_pipe_0 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[1:0];
  _RAND_4 = {16{`RANDOM}};
  data_line_reg = _RAND_4[511:0];
  _RAND_5 = {2{`RANDOM}};
  mem_addr_reg = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  lru_r = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  count = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  Scanf_io_in_valid_REG = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Sram2axi_mulit(
  input         clock,
  input         reset,
  input         io_in_addr_req_valid,
  input  [63:0] io_in_addr_req_bits_addr,
  input         io_in_addr_req_bits_ce,
  input         io_in_addr_req_bits_we,
  output        io_in_rdata_rep_valid,
  output [63:0] io_in_rdata_rep_bits_rdata,
  input  [63:0] io_in_wdata_req_bits_wdata,
  input  [7:0]  io_in_wdata_req_bits_wmask,
  output        io_in_wdata_rep,
  input         io_out_raddr_req_ready,
  output        io_out_raddr_req_valid,
  output [63:0] io_out_raddr_req_bits_addr,
  input         io_out_waddr_req_ready,
  output        io_out_waddr_req_valid,
  output [63:0] io_out_waddr_req_bits_addr,
  output        io_out_rdata_rep_ready,
  input         io_out_rdata_rep_valid,
  input  [63:0] io_out_rdata_rep_bits_rdata,
  output        io_out_wdata_req_valid,
  output [63:0] io_out_wdata_req_bits_wdata,
  output [7:0]  io_out_wdata_req_bits_wmask,
  output        io_out_wb_ready,
  input         io_out_wb_valid,
  input  [1:0]  io_out_wb_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  ar_state; // @[sram2axi.scala 64:25]
  reg  aw_state; // @[sram2axi.scala 65:25]
  wire  _T = ~ar_state; // @[sram2axi.scala 91:19]
  wire  _T_3 = ~io_in_addr_req_bits_we; // @[sram2axi.scala 93:88]
  wire  _GEN_0 = io_in_addr_req_valid & io_out_raddr_req_ready & io_in_addr_req_bits_ce & ~io_in_addr_req_bits_we |
    ar_state; // @[sram2axi.scala 93:112 94:18 64:25]
  wire  _T_7 = ~aw_state; // @[sram2axi.scala 106:20]
  wire  _GEN_4 = io_in_addr_req_valid & io_out_waddr_req_ready & io_in_addr_req_bits_ce & io_in_addr_req_bits_we |
    aw_state; // @[sram2axi.scala 108:112 109:18 65:25]
  wire  _io_out_waddr_req_valid_T_2 = _T_7 & io_in_addr_req_valid & io_in_addr_req_bits_ce; // @[sram2axi.scala 160:75]
  assign io_in_rdata_rep_valid = ar_state & io_out_rdata_rep_valid; // @[sram2axi.scala 154:58]
  assign io_in_rdata_rep_bits_rdata = io_out_rdata_rep_bits_rdata; // @[sram2axi.scala 165:30]
  assign io_in_wdata_rep = io_out_wb_valid & io_out_wb_bits == 2'h0; // @[sram2axi.scala 168:42]
  assign io_out_raddr_req_valid = _T & io_in_addr_req_valid & io_in_addr_req_bits_ce & _T_3; // @[sram2axi.scala 159:101]
  assign io_out_raddr_req_bits_addr = io_in_addr_req_bits_addr; // @[sram2axi.scala 163:30]
  assign io_out_waddr_req_valid = _T_7 & io_in_addr_req_valid & io_in_addr_req_bits_ce & io_in_addr_req_bits_we; // @[sram2axi.scala 160:101]
  assign io_out_waddr_req_bits_addr = io_in_addr_req_bits_addr; // @[sram2axi.scala 164:30]
  assign io_out_rdata_rep_ready = 1'h1; // @[sram2axi.scala 156:26]
  assign io_out_wdata_req_valid = _io_out_waddr_req_valid_T_2 & io_in_addr_req_bits_we; // @[sram2axi.scala 161:101]
  assign io_out_wdata_req_bits_wdata = io_in_wdata_req_bits_wdata; // @[sram2axi.scala 166:31]
  assign io_out_wdata_req_bits_wmask = io_in_wdata_req_bits_wmask; // @[sram2axi.scala 167:31]
  assign io_out_wb_ready = aw_state; // @[sram2axi.scala 157:25]
  always @(posedge clock) begin
    if (reset) begin // @[sram2axi.scala 64:25]
      ar_state <= 1'h0; // @[sram2axi.scala 64:25]
    end else if (~ar_state) begin // @[sram2axi.scala 91:19]
      ar_state <= _GEN_0;
    end else if (ar_state) begin // @[sram2axi.scala 91:19]
      if (io_out_rdata_rep_valid & io_out_rdata_rep_ready) begin // @[sram2axi.scala 100:61]
        ar_state <= 1'h0; // @[sram2axi.scala 101:18]
      end
    end
    if (reset) begin // @[sram2axi.scala 65:25]
      aw_state <= 1'h0; // @[sram2axi.scala 65:25]
    end else if (~aw_state) begin // @[sram2axi.scala 106:20]
      aw_state <= _GEN_4;
    end else if (aw_state) begin // @[sram2axi.scala 106:20]
      if (io_out_wb_valid & io_out_wb_ready) begin // @[sram2axi.scala 115:48]
        aw_state <= 1'h0; // @[sram2axi.scala 116:18]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ar_state = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  aw_state = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AxiArbiter(
  input         clock,
  input         reset,
  output        io_in1_raddr_req_ready,
  input         io_in1_raddr_req_valid,
  input  [63:0] io_in1_raddr_req_bits_addr,
  output        io_in1_waddr_req_ready,
  input         io_in1_waddr_req_valid,
  input  [63:0] io_in1_waddr_req_bits_addr,
  output        io_in1_rdata_rep_valid,
  output [63:0] io_in1_rdata_rep_bits_rdata,
  input         io_in1_wdata_req_valid,
  input  [63:0] io_in1_wdata_req_bits_wdata,
  input  [7:0]  io_in1_wdata_req_bits_wmask,
  input         io_in1_wb_ready,
  output        io_in1_wb_valid,
  output [1:0]  io_in1_wb_bits,
  output        io_in2_raddr_req_ready,
  input         io_in2_raddr_req_valid,
  input  [63:0] io_in2_raddr_req_bits_addr,
  output        io_in2_waddr_req_ready,
  input         io_in2_waddr_req_valid,
  input  [63:0] io_in2_waddr_req_bits_addr,
  output        io_in2_rdata_rep_valid,
  output [63:0] io_in2_rdata_rep_bits_rdata,
  input         io_in2_wdata_req_valid,
  input  [63:0] io_in2_wdata_req_bits_wdata,
  input  [7:0]  io_in2_wdata_req_bits_wmask,
  input         io_in2_wb_ready,
  output        io_in2_wb_valid,
  output [1:0]  io_in2_wb_bits,
  output        io_out_raddr_req_valid,
  output [63:0] io_out_raddr_req_bits_addr,
  output        io_out_waddr_req_valid,
  output [63:0] io_out_waddr_req_bits_addr,
  input         io_out_rdata_rep_valid,
  input  [63:0] io_out_rdata_rep_bits_rdata,
  output        io_out_wdata_req_valid,
  output [63:0] io_out_wdata_req_bits_wdata,
  output [7:0]  io_out_wdata_req_bits_wmask,
  output        io_out_wb_ready,
  input         io_out_wb_valid,
  input  [1:0]  io_out_wb_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  state; // @[AxiArbiter.scala 14:22]
  reg  choose_r; // @[AxiArbiter.scala 15:25]
  wire  _T_1 = ~state; // @[AxiArbiter.scala 17:68]
  wire  _T_5 = (io_in2_raddr_req_valid | io_in2_waddr_req_valid) & _T_1; // @[AxiArbiter.scala 39:65]
  wire  _GEN_0 = (io_in2_raddr_req_valid | io_in2_waddr_req_valid) & _T_1 | choose_r; // @[AxiArbiter.scala 39:83 40:14 15:25]
  wire  _GEN_2 = (io_in2_raddr_req_valid | io_in2_waddr_req_valid) & _T_1 & io_in2_raddr_req_valid; // @[AxiArbiter.scala 39:83 49:28 70:28]
  wire  _GEN_3 = (io_in2_raddr_req_valid | io_in2_waddr_req_valid) & _T_1 & io_in2_waddr_req_valid; // @[AxiArbiter.scala 39:83 50:28 71:28]
  wire  _GEN_4 = (io_in2_raddr_req_valid | io_in2_waddr_req_valid) & _T_1 & io_in2_wdata_req_valid; // @[AxiArbiter.scala 39:83 51:28 72:28]
  wire [63:0] _GEN_6 = (io_in2_raddr_req_valid | io_in2_waddr_req_valid) & _T_1 ? io_in2_raddr_req_bits_addr :
    io_in1_raddr_req_bits_addr; // @[AxiArbiter.scala 39:83 57:27 78:27]
  wire [63:0] _GEN_7 = (io_in2_raddr_req_valid | io_in2_waddr_req_valid) & _T_1 ? io_in2_waddr_req_bits_addr :
    io_in1_waddr_req_bits_addr; // @[AxiArbiter.scala 39:83 58:27 79:27]
  wire [7:0] _GEN_8 = (io_in2_raddr_req_valid | io_in2_waddr_req_valid) & _T_1 ? io_in2_wdata_req_bits_wmask :
    io_in1_wdata_req_bits_wmask; // @[AxiArbiter.scala 39:83 59:27 80:27]
  wire [63:0] _GEN_9 = (io_in2_raddr_req_valid | io_in2_waddr_req_valid) & _T_1 ? io_in2_wdata_req_bits_wdata :
    io_in1_wdata_req_bits_wdata; // @[AxiArbiter.scala 39:83 59:27 80:27]
  wire  _GEN_20 = (io_in1_raddr_req_valid | io_in1_waddr_req_valid) & ~state | _T_5; // @[AxiArbiter.scala 17:77 38:11]
  wire  _GEN_21 = ~choose_r & io_out_rdata_rep_valid; // @[AxiArbiter.scala 85:27 113:30 92:30]
  wire  _GEN_22 = ~choose_r & io_out_wb_valid; // @[AxiArbiter.scala 114:23 85:27 93:23]
  wire  _GEN_23 = ~choose_r ? 1'h0 : io_out_rdata_rep_valid; // @[AxiArbiter.scala 85:27 110:30 95:30]
  wire  _GEN_24 = ~choose_r ? 1'h0 : io_out_wb_valid; // @[AxiArbiter.scala 111:23 85:27 96:23]
  wire  _GEN_26 = ~choose_r ? io_in1_wb_ready : io_in2_wb_ready; // @[AxiArbiter.scala 117:23 85:27 99:23]
  assign io_in1_raddr_req_ready = (io_in1_raddr_req_valid | io_in1_waddr_req_valid) & ~state; // @[AxiArbiter.scala 17:59]
  assign io_in1_waddr_req_ready = (io_in1_raddr_req_valid | io_in1_waddr_req_valid) & ~state; // @[AxiArbiter.scala 17:59]
  assign io_in1_rdata_rep_valid = (io_out_rdata_rep_valid | io_out_wb_valid) & _GEN_21; // @[AxiArbiter.scala 126:28 84:50]
  assign io_in1_rdata_rep_bits_rdata = io_out_rdata_rep_bits_rdata; // @[AxiArbiter.scala 140:25]
  assign io_in1_wb_valid = (io_out_rdata_rep_valid | io_out_wb_valid) & _GEN_22; // @[AxiArbiter.scala 127:21 84:50]
  assign io_in1_wb_bits = io_out_wb_bits; // @[AxiArbiter.scala 141:18]
  assign io_in2_raddr_req_ready = (io_in1_raddr_req_valid | io_in1_waddr_req_valid) & ~state ? 1'h0 : _T_5; // @[AxiArbiter.scala 17:77 31:28]
  assign io_in2_waddr_req_ready = (io_in1_raddr_req_valid | io_in1_waddr_req_valid) & ~state ? 1'h0 : _T_5; // @[AxiArbiter.scala 17:77 31:28]
  assign io_in2_rdata_rep_valid = (io_out_rdata_rep_valid | io_out_wb_valid) & _GEN_23; // @[AxiArbiter.scala 129:28 84:50]
  assign io_in2_rdata_rep_bits_rdata = io_out_rdata_rep_bits_rdata; // @[AxiArbiter.scala 137:25]
  assign io_in2_wb_valid = (io_out_rdata_rep_valid | io_out_wb_valid) & _GEN_24; // @[AxiArbiter.scala 130:21 84:50]
  assign io_in2_wb_bits = io_out_wb_bits; // @[AxiArbiter.scala 138:18]
  assign io_out_raddr_req_valid = (io_in1_raddr_req_valid | io_in1_waddr_req_valid) & ~state ? io_in1_raddr_req_valid :
    _GEN_2; // @[AxiArbiter.scala 17:77 27:28]
  assign io_out_raddr_req_bits_addr = (io_in1_raddr_req_valid | io_in1_waddr_req_valid) & ~state ?
    io_in1_raddr_req_bits_addr : _GEN_6; // @[AxiArbiter.scala 17:77 35:27]
  assign io_out_waddr_req_valid = (io_in1_raddr_req_valid | io_in1_waddr_req_valid) & ~state ? io_in1_waddr_req_valid :
    _GEN_3; // @[AxiArbiter.scala 17:77 28:28]
  assign io_out_waddr_req_bits_addr = (io_in1_raddr_req_valid | io_in1_waddr_req_valid) & ~state ?
    io_in1_waddr_req_bits_addr : _GEN_7; // @[AxiArbiter.scala 17:77 36:27]
  assign io_out_wdata_req_valid = (io_in1_raddr_req_valid | io_in1_waddr_req_valid) & ~state ? io_in1_wdata_req_valid :
    _GEN_4; // @[AxiArbiter.scala 17:77 29:28]
  assign io_out_wdata_req_bits_wdata = (io_in1_raddr_req_valid | io_in1_waddr_req_valid) & ~state ?
    io_in1_wdata_req_bits_wdata : _GEN_9; // @[AxiArbiter.scala 17:77 37:27]
  assign io_out_wdata_req_bits_wmask = (io_in1_raddr_req_valid | io_in1_waddr_req_valid) & ~state ?
    io_in1_wdata_req_bits_wmask : _GEN_8; // @[AxiArbiter.scala 17:77 37:27]
  assign io_out_wb_ready = io_out_rdata_rep_valid | io_out_wb_valid ? _GEN_26 : 1'h1; // @[AxiArbiter.scala 133:21 84:50]
  always @(posedge clock) begin
    if (reset) begin // @[AxiArbiter.scala 14:22]
      state <= 1'h0; // @[AxiArbiter.scala 14:22]
    end else if (io_out_rdata_rep_valid | io_out_wb_valid) begin // @[AxiArbiter.scala 84:50]
      state <= 1'h0;
    end else begin
      state <= _GEN_20;
    end
    if (reset) begin // @[AxiArbiter.scala 15:25]
      choose_r <= 1'h0; // @[AxiArbiter.scala 15:25]
    end else if ((io_in1_raddr_req_valid | io_in1_waddr_req_valid) & ~state) begin // @[AxiArbiter.scala 17:77]
      choose_r <= 1'h0; // @[AxiArbiter.scala 18:14]
    end else begin
      choose_r <= _GEN_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  choose_r = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Cache_1(
  input         clock,
  input         reset,
  input         io_in_addr_req_valid,
  input  [63:0] io_in_addr_req_bits_addr,
  input         io_in_addr_req_bits_we,
  output        io_in_rdata_rep_valid,
  output [63:0] io_in_rdata_rep_bits_rdata,
  input  [63:0] io_in_wdata_req_bits_wdata,
  input  [7:0]  io_in_wdata_req_bits_wmask,
  output        io_in_wdata_rep,
  output        io_out_addr_req_valid,
  output [63:0] io_out_addr_req_bits_addr,
  output        io_out_addr_req_bits_ce,
  output        io_out_addr_req_bits_we,
  input         io_out_rdata_rep_valid,
  input  [63:0] io_out_rdata_rep_bits_rdata,
  output [63:0] io_out_wdata_req_bits_wdata,
  input         io_out_wdata_rep
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [511:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [511:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  Cache_data_clock; // @[Cache.scala 159:26]
  wire  Cache_data_io_in_valid; // @[Cache.scala 159:26]
  wire [63:0] Cache_data_io_in_addr; // @[Cache.scala 159:26]
  wire [63:0] Cache_data_io_write_bus_addr; // @[Cache.scala 159:26]
  wire  Cache_data_io_write_bus_valid; // @[Cache.scala 159:26]
  wire [1:0] Cache_data_io_write_bus_waymask; // @[Cache.scala 159:26]
  wire [511:0] Cache_data_io_write_bus_wdata; // @[Cache.scala 159:26]
  wire  Cache_data_io_out_valid; // @[Cache.scala 159:26]
  wire [52:0] Cache_data_io_out_bits_meat_tag_0; // @[Cache.scala 159:26]
  wire [52:0] Cache_data_io_out_bits_meat_tag_1; // @[Cache.scala 159:26]
  wire  Cache_data_io_out_bits_meat_valid_0; // @[Cache.scala 159:26]
  wire  Cache_data_io_out_bits_meat_valid_1; // @[Cache.scala 159:26]
  wire [511:0] Cache_data_io_out_bits_data_data_0; // @[Cache.scala 159:26]
  wire [511:0] Cache_data_io_out_bits_data_data_1; // @[Cache.scala 159:26]
  wire [52:0] Cache_data_io_out_bits_ctrl_data_tag; // @[Cache.scala 159:26]
  wire [4:0] Cache_data_io_out_bits_ctrl_data_index; // @[Cache.scala 159:26]
  wire [5:0] Cache_data_io_out_bits_ctrl_data_offset; // @[Cache.scala 159:26]
  wire  Scanf_io_in_valid; // @[Cache.scala 160:21]
  wire [52:0] Scanf_io_in_bits_meat_tag_0; // @[Cache.scala 160:21]
  wire [52:0] Scanf_io_in_bits_meat_tag_1; // @[Cache.scala 160:21]
  wire  Scanf_io_in_bits_meat_valid_0; // @[Cache.scala 160:21]
  wire  Scanf_io_in_bits_meat_valid_1; // @[Cache.scala 160:21]
  wire [511:0] Scanf_io_in_bits_data_data_0; // @[Cache.scala 160:21]
  wire [511:0] Scanf_io_in_bits_data_data_1; // @[Cache.scala 160:21]
  wire [52:0] Scanf_io_in_bits_ctrl_data_tag; // @[Cache.scala 160:21]
  wire [4:0] Scanf_io_in_bits_ctrl_data_index; // @[Cache.scala 160:21]
  wire  Scanf_io_out_bits_hit; // @[Cache.scala 160:21]
  wire [511:0] Scanf_io_out_bits_data; // @[Cache.scala 160:21]
  wire [4:0] Scanf_io_out_bits_meta_ctrl_data_index; // @[Cache.scala 160:21]
  wire  Scanf_io_out_bits_hit_way_0; // @[Cache.scala 160:21]
  wire  Scanf_io_out_bits_hit_way_1; // @[Cache.scala 160:21]
  wire [52:0] Scanf_io_out_bits_tag_0; // @[Cache.scala 160:21]
  wire [52:0] Scanf_io_out_bits_tag_1; // @[Cache.scala 160:21]
  reg  lru [0:31]; // @[Cache.scala 173:24]
  wire  lru_lru_w_MPORT_en; // @[Cache.scala 173:24]
  wire [4:0] lru_lru_w_MPORT_addr; // @[Cache.scala 173:24]
  wire  lru_lru_w_MPORT_data; // @[Cache.scala 173:24]
  wire  lru_MPORT_data; // @[Cache.scala 173:24]
  wire [4:0] lru_MPORT_addr; // @[Cache.scala 173:24]
  wire  lru_MPORT_mask; // @[Cache.scala 173:24]
  wire  lru_MPORT_en; // @[Cache.scala 173:24]
  wire  lru_MPORT_1_data; // @[Cache.scala 173:24]
  wire [4:0] lru_MPORT_1_addr; // @[Cache.scala 173:24]
  wire  lru_MPORT_1_mask; // @[Cache.scala 173:24]
  wire  lru_MPORT_1_en; // @[Cache.scala 173:24]
  wire  lru_MPORT_2_data; // @[Cache.scala 173:24]
  wire [4:0] lru_MPORT_2_addr; // @[Cache.scala 173:24]
  wire  lru_MPORT_2_mask; // @[Cache.scala 173:24]
  wire  lru_MPORT_2_en; // @[Cache.scala 173:24]
  wire  lru_MPORT_3_data; // @[Cache.scala 173:24]
  wire [4:0] lru_MPORT_3_addr; // @[Cache.scala 173:24]
  wire  lru_MPORT_3_mask; // @[Cache.scala 173:24]
  wire  lru_MPORT_3_en; // @[Cache.scala 173:24]
  reg  lru_lru_w_MPORT_en_pipe_0;
  reg [4:0] lru_lru_w_MPORT_addr_pipe_0;
  reg  dirt_0 [0:31]; // @[Cache.scala 181:51]
  wire  dirt_0_dirt_w_en; // @[Cache.scala 181:51]
  wire [4:0] dirt_0_dirt_w_addr; // @[Cache.scala 181:51]
  wire  dirt_0_dirt_w_data; // @[Cache.scala 181:51]
  wire  dirt_0_MPORT_4_data; // @[Cache.scala 181:51]
  wire [4:0] dirt_0_MPORT_4_addr; // @[Cache.scala 181:51]
  wire  dirt_0_MPORT_4_mask; // @[Cache.scala 181:51]
  wire  dirt_0_MPORT_4_en; // @[Cache.scala 181:51]
  reg  dirt_0_dirt_w_en_pipe_0;
  reg [4:0] dirt_0_dirt_w_addr_pipe_0;
  reg  dirt_1 [0:31]; // @[Cache.scala 181:51]
  wire  dirt_1_dirt_w_en; // @[Cache.scala 181:51]
  wire [4:0] dirt_1_dirt_w_addr; // @[Cache.scala 181:51]
  wire  dirt_1_dirt_w_data; // @[Cache.scala 181:51]
  wire  dirt_1_MPORT_4_data; // @[Cache.scala 181:51]
  wire [4:0] dirt_1_MPORT_4_addr; // @[Cache.scala 181:51]
  wire  dirt_1_MPORT_4_mask; // @[Cache.scala 181:51]
  wire  dirt_1_MPORT_4_en; // @[Cache.scala 181:51]
  reg  dirt_1_dirt_w_en_pipe_0;
  reg [4:0] dirt_1_dirt_w_addr_pipe_0;
  reg [1:0] state; // @[Cache.scala 163:22]
  reg [511:0] data_line_reg; // @[Cache.scala 165:30]
  reg [63:0] mem_addr_reg; // @[Cache.scala 166:29]
  reg  lru_r; // @[Cache.scala 168:23]
  reg [3:0] count; // @[Cache.scala 176:22]
  wire  s = count == 4'h8; // @[Cache.scala 177:17]
  reg [3:0] count_write; // @[Cache.scala 182:54]
  wire  s_w = count_write == 4'h8; // @[Cache.scala 183:55]
  reg [63:0] mem_write_addr_reg; // @[Cache.scala 185:61]
  reg [511:0] mem_write_data_reg; // @[Cache.scala 186:61]
  wire  _T = 2'h0 == state; // @[Cache.scala 196:16]
  wire  _T_1 = 2'h1 == state; // @[Cache.scala 196:16]
  wire [63:0] _mem_addr_reg_T_2 = {io_in_addr_req_bits_addr[63:6],6'h0}; // @[Cat.scala 31:58]
  wire  lru_w = lru_lru_w_MPORT_data;
  wire [52:0] _GEN_5 = Scanf_io_out_bits_tag_0; // @[Cat.scala 31:{58,58}]
  wire [52:0] _GEN_6 = lru_w ? Scanf_io_out_bits_tag_1 : _GEN_5; // @[Cat.scala 31:{58,58}]
  wire [63:0] _mem_write_addr_reg_T_3 = {_GEN_6,Scanf_io_out_bits_meta_ctrl_data_index,6'h0}; // @[Cat.scala 31:58]
  wire [511:0] _GEN_7 = Cache_data_io_out_bits_data_data_0; // @[Cache.scala 208:{36,36}]
  wire [511:0] _GEN_8 = lru_w ? Cache_data_io_out_bits_data_data_1 : _GEN_7; // @[Cache.scala 208:{36,36}]
  wire  hit_way_0 = Scanf_io_out_bits_hit_way_0; // @[Cache.scala 192:21 357:11]
  wire  hit_way_1 = Scanf_io_out_bits_hit_way_1; // @[Cache.scala 192:21 357:11]
  wire  _GEN_29 = ~Scanf_io_out_bits_hit ? 1'h0 : hit_way_0; // @[Cache.scala 173:24 201:26]
  wire  _GEN_33 = ~Scanf_io_out_bits_hit ? 1'h0 : hit_way_1; // @[Cache.scala 173:24 201:26]
  wire  _T_5 = 2'h2 == state; // @[Cache.scala 196:16]
  wire [3:0] _count_T_1 = count + 4'h1; // @[Cache.scala 229:24]
  wire [63:0] _mem_addr_reg_T_4 = mem_addr_reg + 64'h8; // @[Cache.scala 230:38]
  wire [3:0] _GEN_36 = ~io_out_rdata_rep_valid ? count : _count_T_1; // @[Cache.scala 226:83 227:15 229:15]
  wire [63:0] _GEN_37 = ~io_out_rdata_rep_valid ? mem_addr_reg : _mem_addr_reg_T_4; // @[Cache.scala 166:29 226:83 230:22]
  wire [511:0] _data_line_reg_T_1 = {io_out_rdata_rep_bits_rdata,data_line_reg[511:64]}; // @[Cat.scala 31:58]
  wire [511:0] _GEN_38 = ~s & io_out_rdata_rep_valid ? _data_line_reg_T_1 : data_line_reg; // @[Cache.scala 236:51 237:23 165:30]
  wire  _GEN_46 = lru_r ? 1'h0 : 1'h1; // @[Cache.scala 173:24 240:29]
  wire  _GEN_50 = s & lru_r; // @[Cache.scala 173:24 239:51]
  wire  _GEN_55 = s & _GEN_46; // @[Cache.scala 173:24 239:51]
  wire [3:0] _GEN_57 = s ? 4'h0 : _GEN_36; // @[Cache.scala 239:51 245:14]
  wire  _T_16 = 2'h3 == state; // @[Cache.scala 196:16]
  wire [3:0] _count_write_T_1 = count_write + 4'h1; // @[Cache.scala 252:46]
  wire [63:0] _mem_write_addr_reg_T_5 = mem_write_addr_reg + 64'h8; // @[Cache.scala 253:60]
  wire [511:0] _mem_write_data_reg_T_4 = {64'h0,mem_write_data_reg[511:64]}; // @[Cat.scala 31:58]
  wire [3:0] _GEN_58 = io_out_wdata_rep ? _count_write_T_1 : count_write; // @[Cache.scala 251:35 252:27 182:54]
  wire [63:0] _GEN_59 = io_out_wdata_rep ? _mem_write_addr_reg_T_5 : mem_write_addr_reg; // @[Cache.scala 251:35 253:34 185:61]
  wire [511:0] _GEN_60 = io_out_wdata_rep ? _mem_write_data_reg_T_4 : mem_write_data_reg; // @[Cache.scala 251:35 254:34 186:61]
  wire [3:0] _GEN_61 = s_w ? 4'h0 : _GEN_58; // @[Cache.scala 257:33 258:27]
  wire [3:0] _GEN_62 = 2'h3 == state ? _GEN_61 : count_write; // @[Cache.scala 196:16 182:54]
  wire [63:0] _GEN_63 = 2'h3 == state ? _GEN_59 : mem_write_addr_reg; // @[Cache.scala 196:16 185:61]
  wire [511:0] _GEN_64 = 2'h3 == state ? _GEN_60 : mem_write_data_reg; // @[Cache.scala 196:16 186:61]
  wire  _GEN_91 = 2'h1 == state & _GEN_29; // @[Cache.scala 196:16 173:24]
  wire  _GEN_95 = 2'h1 == state & _GEN_33; // @[Cache.scala 196:16 173:24]
  wire  _GEN_102 = 2'h1 == state ? 1'h0 : 2'h2 == state & _GEN_50; // @[Cache.scala 196:16 173:24]
  wire  _GEN_107 = 2'h1 == state ? 1'h0 : 2'h2 == state & _GEN_55; // @[Cache.scala 196:16 173:24]
  wire [63:0] _GEN_138 = 3'h7 == io_in_addr_req_bits_addr[5:3] ? Scanf_io_out_bits_data[511:448] : 64'h0; // @[Cache.scala 266:115 296:16]
  wire [63:0] _GEN_139 = 3'h7 == io_in_addr_req_bits_addr[5:3] ? data_line_reg[511:448] : 64'h0; // @[Cache.scala 266:115 297:16]
  wire [63:0] _GEN_140 = 3'h6 == io_in_addr_req_bits_addr[5:3] ? Scanf_io_out_bits_data[447:384] : _GEN_138; // @[Cache.scala 266:115 292:16]
  wire [63:0] _GEN_141 = 3'h6 == io_in_addr_req_bits_addr[5:3] ? data_line_reg[447:384] : _GEN_139; // @[Cache.scala 266:115 293:16]
  wire [63:0] _GEN_142 = 3'h5 == io_in_addr_req_bits_addr[5:3] ? Scanf_io_out_bits_data[383:320] : _GEN_140; // @[Cache.scala 266:115 288:16]
  wire [63:0] _GEN_143 = 3'h5 == io_in_addr_req_bits_addr[5:3] ? data_line_reg[383:320] : _GEN_141; // @[Cache.scala 266:115 289:16]
  wire [63:0] _GEN_144 = 3'h4 == io_in_addr_req_bits_addr[5:3] ? Scanf_io_out_bits_data[319:256] : _GEN_142; // @[Cache.scala 266:115 284:16]
  wire [63:0] _GEN_145 = 3'h4 == io_in_addr_req_bits_addr[5:3] ? data_line_reg[319:256] : _GEN_143; // @[Cache.scala 266:115 285:16]
  wire [63:0] _GEN_146 = 3'h3 == io_in_addr_req_bits_addr[5:3] ? Scanf_io_out_bits_data[255:192] : _GEN_144; // @[Cache.scala 266:115 280:16]
  wire [63:0] _GEN_147 = 3'h3 == io_in_addr_req_bits_addr[5:3] ? data_line_reg[255:192] : _GEN_145; // @[Cache.scala 266:115 281:16]
  wire [63:0] _GEN_148 = 3'h2 == io_in_addr_req_bits_addr[5:3] ? Scanf_io_out_bits_data[191:128] : _GEN_146; // @[Cache.scala 266:115 276:16]
  wire [63:0] _GEN_149 = 3'h2 == io_in_addr_req_bits_addr[5:3] ? data_line_reg[191:128] : _GEN_147; // @[Cache.scala 266:115 277:16]
  wire [63:0] _GEN_150 = 3'h1 == io_in_addr_req_bits_addr[5:3] ? Scanf_io_out_bits_data[127:64] : _GEN_148; // @[Cache.scala 266:115 272:16]
  wire [63:0] _GEN_151 = 3'h1 == io_in_addr_req_bits_addr[5:3] ? data_line_reg[127:64] : _GEN_149; // @[Cache.scala 266:115 273:16]
  wire [63:0] hit_data = 3'h0 == io_in_addr_req_bits_addr[5:3] ? Scanf_io_out_bits_data[63:0] : _GEN_150; // @[Cache.scala 266:115 268:16]
  wire [63:0] mem_data = 3'h0 == io_in_addr_req_bits_addr[5:3] ? data_line_reg[63:0] : _GEN_151; // @[Cache.scala 266:115 269:16]
  wire  _GEN_156 = lru_w ? dirt_1_dirt_w_data : dirt_0_dirt_w_data; // @[Cache.scala 314:{36,36}]
  wire [1:0] _GEN_157 = _GEN_156 ? 2'h3 : 2'h2; // @[Cache.scala 314:44 315:21 317:21]
  wire [1:0] _GEN_159 = s ? 2'h0 : state; // @[Cache.scala 327:52 328:17 163:22]
  wire [1:0] _GEN_160 = s_w ? 2'h2 : state; // @[Cache.scala 334:34 335:17 163:22]
  wire [1:0] _GEN_161 = _T_16 ? _GEN_160 : state; // @[Cache.scala 301:16 163:22]
  wire  _io_in_rdata_rep_bits_rdata_T = state == 2'h1; // @[Cache.scala 345:44]
  wire  _io_in_rdata_rep_bits_rdata_T_1 = state == 2'h1 & Scanf_io_out_bits_hit; // @[Cache.scala 345:54]
  reg  Scanf_io_in_valid_REG; // @[Cache.scala 352:31]
  wire  _io_out_addr_req_valid_T = state == 2'h2; // @[Cache.scala 364:40]
  wire  _io_out_addr_req_valid_T_1 = state == 2'h3; // @[Cache.scala 364:58]
  wire  _io_out_addr_req_bits_ce_T_2 = ~s_w; // @[Cache.scala 365:79]
  wire  _io_in_rdata_rep_valid_T_4 = _io_out_addr_req_valid_T & s; // @[Cache.scala 381:75]
  wire  _io_in_rdata_rep_valid_T_5 = _io_in_rdata_rep_bits_rdata_T_1 | _io_out_addr_req_valid_T & s; // @[Cache.scala 381:57]
  wire [7:0] _wmaskextend_T_2 = io_in_addr_req_bits_we ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_3 = io_in_wdata_req_bits_wmask & _wmaskextend_T_2; // @[Cache.scala 384:38]
  wire  _wmaskextend_Genmask_T = Cache_data_io_out_bits_ctrl_data_offset[5:3] == 3'h0; // @[util.scala 55:15]
  wire [63:0] _wmaskextend_Genmask_T_2 = {56'h0,_wmaskextend_T_3}; // @[Cat.scala 31:58]
  wire  _wmaskextend_Genmask_T_3 = Cache_data_io_out_bits_ctrl_data_offset[5:3] == 3'h1; // @[util.scala 56:15]
  wire [63:0] _wmaskextend_Genmask_T_6 = {48'h0,_wmaskextend_T_3,8'h0}; // @[Cat.scala 31:58]
  wire  _wmaskextend_Genmask_T_7 = Cache_data_io_out_bits_ctrl_data_offset[5:3] == 3'h2; // @[util.scala 57:15]
  wire [63:0] _wmaskextend_Genmask_T_10 = {40'h0,_wmaskextend_T_3,16'h0}; // @[Cat.scala 31:58]
  wire  _wmaskextend_Genmask_T_11 = Cache_data_io_out_bits_ctrl_data_offset[5:3] == 3'h3; // @[util.scala 58:15]
  wire [63:0] _wmaskextend_Genmask_T_14 = {32'h0,_wmaskextend_T_3,24'h0}; // @[Cat.scala 31:58]
  wire  _wmaskextend_Genmask_T_15 = Cache_data_io_out_bits_ctrl_data_offset[5:3] == 3'h4; // @[util.scala 59:15]
  wire [63:0] _wmaskextend_Genmask_T_18 = {24'h0,_wmaskextend_T_3,32'h0}; // @[Cat.scala 31:58]
  wire  _wmaskextend_Genmask_T_19 = Cache_data_io_out_bits_ctrl_data_offset[5:3] == 3'h5; // @[util.scala 60:15]
  wire [63:0] _wmaskextend_Genmask_T_22 = {16'h0,_wmaskextend_T_3,40'h0}; // @[Cat.scala 31:58]
  wire  _wmaskextend_Genmask_T_23 = Cache_data_io_out_bits_ctrl_data_offset[5:3] == 3'h6; // @[util.scala 61:15]
  wire [63:0] _wmaskextend_Genmask_T_26 = {8'h0,_wmaskextend_T_3,48'h0}; // @[Cat.scala 31:58]
  wire  _wmaskextend_Genmask_T_27 = Cache_data_io_out_bits_ctrl_data_offset[5:3] == 3'h7; // @[util.scala 62:15]
  wire [63:0] _wmaskextend_Genmask_T_29 = {_wmaskextend_T_3,56'h0}; // @[Cat.scala 31:58]
  wire [63:0] _wmaskextend_Genmask_T_30 = _wmaskextend_Genmask_T_27 ? _wmaskextend_Genmask_T_29 : 64'h0; // @[Mux.scala 101:16]
  wire [63:0] _wmaskextend_Genmask_T_31 = _wmaskextend_Genmask_T_23 ? _wmaskextend_Genmask_T_26 :
    _wmaskextend_Genmask_T_30; // @[Mux.scala 101:16]
  wire [63:0] _wmaskextend_Genmask_T_32 = _wmaskextend_Genmask_T_19 ? _wmaskextend_Genmask_T_22 :
    _wmaskextend_Genmask_T_31; // @[Mux.scala 101:16]
  wire [63:0] _wmaskextend_Genmask_T_33 = _wmaskextend_Genmask_T_15 ? _wmaskextend_Genmask_T_18 :
    _wmaskextend_Genmask_T_32; // @[Mux.scala 101:16]
  wire [63:0] _wmaskextend_Genmask_T_34 = _wmaskextend_Genmask_T_11 ? _wmaskextend_Genmask_T_14 :
    _wmaskextend_Genmask_T_33; // @[Mux.scala 101:16]
  wire [63:0] _wmaskextend_Genmask_T_35 = _wmaskextend_Genmask_T_7 ? _wmaskextend_Genmask_T_10 :
    _wmaskextend_Genmask_T_34; // @[Mux.scala 101:16]
  wire [63:0] _wmaskextend_Genmask_T_36 = _wmaskextend_Genmask_T_3 ? _wmaskextend_Genmask_T_6 :
    _wmaskextend_Genmask_T_35; // @[Mux.scala 101:16]
  wire [63:0] wmaskextend_Genmask = _wmaskextend_Genmask_T ? _wmaskextend_Genmask_T_2 : _wmaskextend_Genmask_T_36; // @[Mux.scala 101:16]
  wire [7:0] _wmaskextend_T_69 = wmaskextend_Genmask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_71 = wmaskextend_Genmask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_73 = wmaskextend_Genmask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_75 = wmaskextend_Genmask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_77 = wmaskextend_Genmask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_79 = wmaskextend_Genmask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_81 = wmaskextend_Genmask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_83 = wmaskextend_Genmask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_85 = wmaskextend_Genmask[8] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_87 = wmaskextend_Genmask[9] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_89 = wmaskextend_Genmask[10] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_91 = wmaskextend_Genmask[11] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_93 = wmaskextend_Genmask[12] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_95 = wmaskextend_Genmask[13] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_97 = wmaskextend_Genmask[14] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_99 = wmaskextend_Genmask[15] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_101 = wmaskextend_Genmask[16] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_103 = wmaskextend_Genmask[17] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_105 = wmaskextend_Genmask[18] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_107 = wmaskextend_Genmask[19] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_109 = wmaskextend_Genmask[20] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_111 = wmaskextend_Genmask[21] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_113 = wmaskextend_Genmask[22] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_115 = wmaskextend_Genmask[23] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_117 = wmaskextend_Genmask[24] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_119 = wmaskextend_Genmask[25] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_121 = wmaskextend_Genmask[26] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_123 = wmaskextend_Genmask[27] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_125 = wmaskextend_Genmask[28] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_127 = wmaskextend_Genmask[29] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_129 = wmaskextend_Genmask[30] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_131 = wmaskextend_Genmask[31] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_133 = wmaskextend_Genmask[32] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_135 = wmaskextend_Genmask[33] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_137 = wmaskextend_Genmask[34] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_139 = wmaskextend_Genmask[35] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_141 = wmaskextend_Genmask[36] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_143 = wmaskextend_Genmask[37] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_145 = wmaskextend_Genmask[38] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_147 = wmaskextend_Genmask[39] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_149 = wmaskextend_Genmask[40] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_151 = wmaskextend_Genmask[41] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_153 = wmaskextend_Genmask[42] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_155 = wmaskextend_Genmask[43] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_157 = wmaskextend_Genmask[44] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_159 = wmaskextend_Genmask[45] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_161 = wmaskextend_Genmask[46] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_163 = wmaskextend_Genmask[47] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_165 = wmaskextend_Genmask[48] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_167 = wmaskextend_Genmask[49] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_169 = wmaskextend_Genmask[50] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_171 = wmaskextend_Genmask[51] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_173 = wmaskextend_Genmask[52] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_175 = wmaskextend_Genmask[53] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_177 = wmaskextend_Genmask[54] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_179 = wmaskextend_Genmask[55] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_181 = wmaskextend_Genmask[56] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_183 = wmaskextend_Genmask[57] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_185 = wmaskextend_Genmask[58] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_187 = wmaskextend_Genmask[59] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_189 = wmaskextend_Genmask[60] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_191 = wmaskextend_Genmask[61] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_193 = wmaskextend_Genmask[62] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wmaskextend_T_195 = wmaskextend_Genmask[63] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [63:0] wmaskextend_lo_lo_lo = {_wmaskextend_T_83,_wmaskextend_T_81,_wmaskextend_T_79,_wmaskextend_T_77,
    _wmaskextend_T_75,_wmaskextend_T_73,_wmaskextend_T_71,_wmaskextend_T_69}; // @[Cat.scala 31:58]
  wire [127:0] wmaskextend_lo_lo = {_wmaskextend_T_99,_wmaskextend_T_97,_wmaskextend_T_95,_wmaskextend_T_93,
    _wmaskextend_T_91,_wmaskextend_T_89,_wmaskextend_T_87,_wmaskextend_T_85,wmaskextend_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [63:0] wmaskextend_lo_hi_lo = {_wmaskextend_T_115,_wmaskextend_T_113,_wmaskextend_T_111,_wmaskextend_T_109,
    _wmaskextend_T_107,_wmaskextend_T_105,_wmaskextend_T_103,_wmaskextend_T_101}; // @[Cat.scala 31:58]
  wire [255:0] wmaskextend_lo = {_wmaskextend_T_131,_wmaskextend_T_129,_wmaskextend_T_127,_wmaskextend_T_125,
    _wmaskextend_T_123,_wmaskextend_T_121,_wmaskextend_T_119,_wmaskextend_T_117,wmaskextend_lo_hi_lo,wmaskextend_lo_lo}; // @[Cat.scala 31:58]
  wire [63:0] wmaskextend_hi_lo_lo = {_wmaskextend_T_147,_wmaskextend_T_145,_wmaskextend_T_143,_wmaskextend_T_141,
    _wmaskextend_T_139,_wmaskextend_T_137,_wmaskextend_T_135,_wmaskextend_T_133}; // @[Cat.scala 31:58]
  wire [127:0] wmaskextend_hi_lo = {_wmaskextend_T_163,_wmaskextend_T_161,_wmaskextend_T_159,_wmaskextend_T_157,
    _wmaskextend_T_155,_wmaskextend_T_153,_wmaskextend_T_151,_wmaskextend_T_149,wmaskextend_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [63:0] wmaskextend_hi_hi_lo = {_wmaskextend_T_179,_wmaskextend_T_177,_wmaskextend_T_175,_wmaskextend_T_173,
    _wmaskextend_T_171,_wmaskextend_T_169,_wmaskextend_T_167,_wmaskextend_T_165}; // @[Cat.scala 31:58]
  wire [255:0] wmaskextend_hi = {_wmaskextend_T_195,_wmaskextend_T_193,_wmaskextend_T_191,_wmaskextend_T_189,
    _wmaskextend_T_187,_wmaskextend_T_185,_wmaskextend_T_183,_wmaskextend_T_181,wmaskextend_hi_hi_lo,wmaskextend_hi_lo}; // @[Cat.scala 31:58]
  wire [511:0] wmaskextend = {wmaskextend_hi,wmaskextend_lo}; // @[Cat.scala 31:58]
  wire [511:0] wdata_extend = {io_in_wdata_req_bits_wdata,io_in_wdata_req_bits_wdata,io_in_wdata_req_bits_wdata,
    io_in_wdata_req_bits_wdata,io_in_wdata_req_bits_wdata,io_in_wdata_req_bits_wdata,io_in_wdata_req_bits_wdata,
    io_in_wdata_req_bits_wdata}; // @[Cat.scala 31:58]
  wire [511:0] _wdata_T_3 = ~wmaskextend; // @[util.scala 38:17]
  wire [511:0] _wdata_T_5 = data_line_reg & _wdata_T_3; // @[util.scala 38:14]
  wire [511:0] _wdata_T_6 = wdata_extend & wmaskextend; // @[util.scala 38:55]
  wire [511:0] _wdata_T_7 = _wdata_T_5 | _wdata_T_6; // @[util.scala 38:44]
  wire [511:0] _wdata_T_10 = Scanf_io_out_bits_data & _wdata_T_3; // @[util.scala 38:14]
  wire [511:0] _wdata_T_12 = _wdata_T_10 | _wdata_T_6; // @[util.scala 38:44]
  wire  _Cache_data_io_write_bus_valid_T_2 = _io_in_rdata_rep_bits_rdata_T & io_in_addr_req_bits_we &
    Scanf_io_out_bits_hit; // @[Cache.scala 397:91]
  wire [1:0] _waymask_T_3 = {hit_way_1,hit_way_0}; // @[Cache.scala 410:80]
  wire [1:0] _waymask_T_5 = lru_r ? 2'h2 : 2'h1; // @[Cache.scala 410:90]
  wire [1:0] waymask = _io_in_rdata_rep_bits_rdata_T_1 & io_in_addr_req_bits_we ? _waymask_T_3 : _waymask_T_5; // @[Cache.scala 410:22]
  Cache_Data Cache_data ( // @[Cache.scala 159:26]
    .clock(Cache_data_clock),
    .io_in_valid(Cache_data_io_in_valid),
    .io_in_addr(Cache_data_io_in_addr),
    .io_write_bus_addr(Cache_data_io_write_bus_addr),
    .io_write_bus_valid(Cache_data_io_write_bus_valid),
    .io_write_bus_waymask(Cache_data_io_write_bus_waymask),
    .io_write_bus_wdata(Cache_data_io_write_bus_wdata),
    .io_out_valid(Cache_data_io_out_valid),
    .io_out_bits_meat_tag_0(Cache_data_io_out_bits_meat_tag_0),
    .io_out_bits_meat_tag_1(Cache_data_io_out_bits_meat_tag_1),
    .io_out_bits_meat_valid_0(Cache_data_io_out_bits_meat_valid_0),
    .io_out_bits_meat_valid_1(Cache_data_io_out_bits_meat_valid_1),
    .io_out_bits_data_data_0(Cache_data_io_out_bits_data_data_0),
    .io_out_bits_data_data_1(Cache_data_io_out_bits_data_data_1),
    .io_out_bits_ctrl_data_tag(Cache_data_io_out_bits_ctrl_data_tag),
    .io_out_bits_ctrl_data_index(Cache_data_io_out_bits_ctrl_data_index),
    .io_out_bits_ctrl_data_offset(Cache_data_io_out_bits_ctrl_data_offset)
  );
  Scanf_data Scanf ( // @[Cache.scala 160:21]
    .io_in_valid(Scanf_io_in_valid),
    .io_in_bits_meat_tag_0(Scanf_io_in_bits_meat_tag_0),
    .io_in_bits_meat_tag_1(Scanf_io_in_bits_meat_tag_1),
    .io_in_bits_meat_valid_0(Scanf_io_in_bits_meat_valid_0),
    .io_in_bits_meat_valid_1(Scanf_io_in_bits_meat_valid_1),
    .io_in_bits_data_data_0(Scanf_io_in_bits_data_data_0),
    .io_in_bits_data_data_1(Scanf_io_in_bits_data_data_1),
    .io_in_bits_ctrl_data_tag(Scanf_io_in_bits_ctrl_data_tag),
    .io_in_bits_ctrl_data_index(Scanf_io_in_bits_ctrl_data_index),
    .io_out_bits_hit(Scanf_io_out_bits_hit),
    .io_out_bits_data(Scanf_io_out_bits_data),
    .io_out_bits_meta_ctrl_data_index(Scanf_io_out_bits_meta_ctrl_data_index),
    .io_out_bits_hit_way_0(Scanf_io_out_bits_hit_way_0),
    .io_out_bits_hit_way_1(Scanf_io_out_bits_hit_way_1),
    .io_out_bits_tag_0(Scanf_io_out_bits_tag_0),
    .io_out_bits_tag_1(Scanf_io_out_bits_tag_1)
  );
  assign lru_lru_w_MPORT_en = lru_lru_w_MPORT_en_pipe_0;
  assign lru_lru_w_MPORT_addr = lru_lru_w_MPORT_addr_pipe_0;
  assign lru_lru_w_MPORT_data = lru[lru_lru_w_MPORT_addr]; // @[Cache.scala 173:24]
  assign lru_MPORT_data = 1'h1;
  assign lru_MPORT_addr = Cache_data_io_out_bits_ctrl_data_index;
  assign lru_MPORT_mask = 1'h1;
  assign lru_MPORT_en = _T ? 1'h0 : _GEN_91;
  assign lru_MPORT_1_data = 1'h0;
  assign lru_MPORT_1_addr = Cache_data_io_out_bits_ctrl_data_index;
  assign lru_MPORT_1_mask = 1'h1;
  assign lru_MPORT_1_en = _T ? 1'h0 : _GEN_95;
  assign lru_MPORT_2_data = 1'h0;
  assign lru_MPORT_2_addr = Cache_data_io_out_bits_ctrl_data_index;
  assign lru_MPORT_2_mask = 1'h1;
  assign lru_MPORT_2_en = _T ? 1'h0 : _GEN_102;
  assign lru_MPORT_3_data = 1'h1;
  assign lru_MPORT_3_addr = Cache_data_io_out_bits_ctrl_data_index;
  assign lru_MPORT_3_mask = 1'h1;
  assign lru_MPORT_3_en = _T ? 1'h0 : _GEN_107;
  assign dirt_0_dirt_w_en = dirt_0_dirt_w_en_pipe_0;
  assign dirt_0_dirt_w_addr = dirt_0_dirt_w_addr_pipe_0;
  assign dirt_0_dirt_w_data = dirt_0[dirt_0_dirt_w_addr]; // @[Cache.scala 181:51]
  assign dirt_0_MPORT_4_data = 1'h1;
  assign dirt_0_MPORT_4_addr = Cache_data_io_out_bits_ctrl_data_index;
  assign dirt_0_MPORT_4_mask = waymask[0];
  assign dirt_0_MPORT_4_en = io_in_addr_req_bits_we & _io_in_rdata_rep_valid_T_5;
  assign dirt_1_dirt_w_en = dirt_1_dirt_w_en_pipe_0;
  assign dirt_1_dirt_w_addr = dirt_1_dirt_w_addr_pipe_0;
  assign dirt_1_dirt_w_data = dirt_1[dirt_1_dirt_w_addr]; // @[Cache.scala 181:51]
  assign dirt_1_MPORT_4_data = 1'h1;
  assign dirt_1_MPORT_4_addr = Cache_data_io_out_bits_ctrl_data_index;
  assign dirt_1_MPORT_4_mask = waymask[1];
  assign dirt_1_MPORT_4_en = io_in_addr_req_bits_we & _io_in_rdata_rep_valid_T_5;
  assign io_in_rdata_rep_valid = (_io_in_rdata_rep_bits_rdata_T_1 | _io_out_addr_req_valid_T & s) & ~
    io_in_addr_req_bits_we; // @[Cache.scala 381:108]
  assign io_in_rdata_rep_bits_rdata = state == 2'h1 & Scanf_io_out_bits_hit ? hit_data : mem_data; // @[Cache.scala 345:36]
  assign io_in_wdata_rep = _Cache_data_io_write_bus_valid_T_2 | _io_in_rdata_rep_valid_T_4 & io_in_addr_req_bits_we; // @[Cache.scala 402:83]
  assign io_out_addr_req_valid = state == 2'h2 | state == 2'h3; // @[Cache.scala 364:49]
  assign io_out_addr_req_bits_addr = _io_out_addr_req_valid_T_1 ? mem_write_addr_reg : mem_addr_reg; // @[Cache.scala 366:37]
  assign io_out_addr_req_bits_ce = _io_out_addr_req_valid_T | _io_out_addr_req_valid_T_1 & ~s_w; // @[Cache.scala 365:51]
  assign io_out_addr_req_bits_we = _io_out_addr_req_valid_T_1 & _io_out_addr_req_bits_ce_T_2; // @[Cache.scala 367:57]
  assign io_out_wdata_req_bits_wdata = mem_write_data_reg[63:0]; // @[Cache.scala 368:62]
  assign Cache_data_clock = clock;
  assign Cache_data_io_in_valid = io_in_addr_req_valid & state == 2'h0; // @[Cache.scala 350:54]
  assign Cache_data_io_in_addr = io_in_addr_req_bits_addr; // @[Cache.scala 351:25]
  assign Cache_data_io_write_bus_addr = _io_in_rdata_rep_valid_T_4 | _Cache_data_io_write_bus_valid_T_2 ?
    io_in_addr_req_bits_addr : 64'h0; // @[Cache.scala 398:40]
  assign Cache_data_io_write_bus_valid = s | _io_in_rdata_rep_bits_rdata_T & io_in_addr_req_bits_we &
    Scanf_io_out_bits_hit; // @[Cache.scala 397:45]
  assign Cache_data_io_write_bus_waymask = _io_in_rdata_rep_bits_rdata_T_1 & io_in_addr_req_bits_we ? _waymask_T_3 :
    _waymask_T_5; // @[Cache.scala 410:22]
  assign Cache_data_io_write_bus_wdata = _io_in_rdata_rep_valid_T_4 ? _wdata_T_7 : _wdata_T_12; // @[Cache.scala 388:20]
  assign Scanf_io_in_valid = Scanf_io_in_valid_REG; // @[Cache.scala 352:21]
  assign Scanf_io_in_bits_meat_tag_0 = Cache_data_io_out_bits_meat_tag_0; // @[Cache.scala 353:25]
  assign Scanf_io_in_bits_meat_tag_1 = Cache_data_io_out_bits_meat_tag_1; // @[Cache.scala 353:25]
  assign Scanf_io_in_bits_meat_valid_0 = Cache_data_io_out_bits_meat_valid_0; // @[Cache.scala 353:25]
  assign Scanf_io_in_bits_meat_valid_1 = Cache_data_io_out_bits_meat_valid_1; // @[Cache.scala 353:25]
  assign Scanf_io_in_bits_data_data_0 = Cache_data_io_out_bits_data_data_0; // @[Cache.scala 354:25]
  assign Scanf_io_in_bits_data_data_1 = Cache_data_io_out_bits_data_data_1; // @[Cache.scala 354:25]
  assign Scanf_io_in_bits_ctrl_data_tag = Cache_data_io_out_bits_ctrl_data_tag; // @[Cache.scala 355:30]
  assign Scanf_io_in_bits_ctrl_data_index = Cache_data_io_out_bits_ctrl_data_index; // @[Cache.scala 355:30]
  always @(posedge clock) begin
    if (lru_MPORT_en & lru_MPORT_mask) begin
      lru[lru_MPORT_addr] <= lru_MPORT_data; // @[Cache.scala 173:24]
    end
    if (lru_MPORT_1_en & lru_MPORT_1_mask) begin
      lru[lru_MPORT_1_addr] <= lru_MPORT_1_data; // @[Cache.scala 173:24]
    end
    if (lru_MPORT_2_en & lru_MPORT_2_mask) begin
      lru[lru_MPORT_2_addr] <= lru_MPORT_2_data; // @[Cache.scala 173:24]
    end
    if (lru_MPORT_3_en & lru_MPORT_3_mask) begin
      lru[lru_MPORT_3_addr] <= lru_MPORT_3_data; // @[Cache.scala 173:24]
    end
    lru_lru_w_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      lru_lru_w_MPORT_addr_pipe_0 <= Cache_data_io_out_bits_ctrl_data_index;
    end
    if (dirt_0_MPORT_4_en & dirt_0_MPORT_4_mask) begin
      dirt_0[dirt_0_MPORT_4_addr] <= dirt_0_MPORT_4_data; // @[Cache.scala 181:51]
    end
    dirt_0_dirt_w_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dirt_0_dirt_w_addr_pipe_0 <= Cache_data_io_out_bits_ctrl_data_index;
    end
    if (dirt_1_MPORT_4_en & dirt_1_MPORT_4_mask) begin
      dirt_1[dirt_1_MPORT_4_addr] <= dirt_1_MPORT_4_data; // @[Cache.scala 181:51]
    end
    dirt_1_dirt_w_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      dirt_1_dirt_w_addr_pipe_0 <= Cache_data_io_out_bits_ctrl_data_index;
    end
    if (reset) begin // @[Cache.scala 163:22]
      state <= 2'h0; // @[Cache.scala 163:22]
    end else if (_T) begin // @[Cache.scala 301:16]
      if (io_in_addr_req_valid) begin // @[Cache.scala 303:33]
        state <= 2'h1; // @[Cache.scala 304:15]
      end else begin
        state <= 2'h0; // @[Cache.scala 306:15]
      end
    end else if (_T_1) begin // @[Cache.scala 301:16]
      if (Scanf_io_out_bits_hit) begin // @[Cache.scala 310:26]
        state <= 2'h0; // @[Cache.scala 311:17]
      end else begin
        state <= _GEN_157;
      end
    end else if (_T_5) begin // @[Cache.scala 301:16]
      state <= _GEN_159;
    end else begin
      state <= _GEN_161;
    end
    if (reset) begin // @[Cache.scala 165:30]
      data_line_reg <= 512'h0; // @[Cache.scala 165:30]
    end else if (!(2'h0 == state)) begin // @[Cache.scala 196:16]
      if (!(2'h1 == state)) begin // @[Cache.scala 196:16]
        if (2'h2 == state) begin // @[Cache.scala 196:16]
          data_line_reg <= _GEN_38;
        end
      end
    end
    if (reset) begin // @[Cache.scala 166:29]
      mem_addr_reg <= 64'h0; // @[Cache.scala 166:29]
    end else if (!(2'h0 == state)) begin // @[Cache.scala 196:16]
      if (2'h1 == state) begin // @[Cache.scala 196:16]
        if (~Scanf_io_out_bits_hit) begin // @[Cache.scala 201:26]
          mem_addr_reg <= _mem_addr_reg_T_2; // @[Cache.scala 202:24]
        end
      end else if (2'h2 == state) begin // @[Cache.scala 196:16]
        mem_addr_reg <= _GEN_37;
      end
    end
    if (reset) begin // @[Cache.scala 168:23]
      lru_r <= 1'h0; // @[Cache.scala 168:23]
    end else if (!(2'h0 == state)) begin // @[Cache.scala 196:16]
      if (2'h1 == state) begin // @[Cache.scala 196:16]
        if (~Scanf_io_out_bits_hit) begin // @[Cache.scala 201:26]
          lru_r <= lru_w; // @[Cache.scala 203:17]
        end
      end
    end
    if (reset) begin // @[Cache.scala 176:22]
      count <= 4'h0; // @[Cache.scala 176:22]
    end else if (2'h0 == state) begin // @[Cache.scala 196:16]
      count <= 4'h0; // @[Cache.scala 198:13]
    end else if (!(2'h1 == state)) begin // @[Cache.scala 196:16]
      if (2'h2 == state) begin // @[Cache.scala 196:16]
        count <= _GEN_57;
      end
    end
    if (reset) begin // @[Cache.scala 182:54]
      count_write <= 4'h0; // @[Cache.scala 182:54]
    end else if (!(2'h0 == state)) begin // @[Cache.scala 196:16]
      if (2'h1 == state) begin // @[Cache.scala 196:16]
        if (~Scanf_io_out_bits_hit) begin // @[Cache.scala 201:26]
          count_write <= 4'h0; // @[Cache.scala 206:29]
        end
      end else if (!(2'h2 == state)) begin // @[Cache.scala 196:16]
        count_write <= _GEN_62;
      end
    end
    if (reset) begin // @[Cache.scala 185:61]
      mem_write_addr_reg <= 64'h0; // @[Cache.scala 185:61]
    end else if (!(2'h0 == state)) begin // @[Cache.scala 196:16]
      if (2'h1 == state) begin // @[Cache.scala 196:16]
        if (~Scanf_io_out_bits_hit) begin // @[Cache.scala 201:26]
          mem_write_addr_reg <= _mem_write_addr_reg_T_3; // @[Cache.scala 207:36]
        end
      end else if (!(2'h2 == state)) begin // @[Cache.scala 196:16]
        mem_write_addr_reg <= _GEN_63;
      end
    end
    if (reset) begin // @[Cache.scala 186:61]
      mem_write_data_reg <= 512'h0; // @[Cache.scala 186:61]
    end else if (!(2'h0 == state)) begin // @[Cache.scala 196:16]
      if (2'h1 == state) begin // @[Cache.scala 196:16]
        if (~Scanf_io_out_bits_hit) begin // @[Cache.scala 201:26]
          mem_write_data_reg <= _GEN_8; // @[Cache.scala 208:36]
        end
      end else if (!(2'h2 == state)) begin // @[Cache.scala 196:16]
        mem_write_data_reg <= _GEN_64;
      end
    end
    Scanf_io_in_valid_REG <= Cache_data_io_out_valid; // @[Cache.scala 352:31]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    lru[initvar] = _RAND_0[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    dirt_0[initvar] = _RAND_3[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    dirt_1[initvar] = _RAND_6[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  lru_lru_w_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  lru_lru_w_MPORT_addr_pipe_0 = _RAND_2[4:0];
  _RAND_4 = {1{`RANDOM}};
  dirt_0_dirt_w_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  dirt_0_dirt_w_addr_pipe_0 = _RAND_5[4:0];
  _RAND_7 = {1{`RANDOM}};
  dirt_1_dirt_w_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  dirt_1_dirt_w_addr_pipe_0 = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  state = _RAND_9[1:0];
  _RAND_10 = {16{`RANDOM}};
  data_line_reg = _RAND_10[511:0];
  _RAND_11 = {2{`RANDOM}};
  mem_addr_reg = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  lru_r = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  count = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  count_write = _RAND_14[3:0];
  _RAND_15 = {2{`RANDOM}};
  mem_write_addr_reg = _RAND_15[63:0];
  _RAND_16 = {16{`RANDOM}};
  mem_write_data_reg = _RAND_16[511:0];
  _RAND_17 = {1{`RANDOM}};
  Scanf_io_in_valid_REG = _RAND_17[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MMIO(
  input         clock,
  input         reset,
  input         io_in_addr_req_valid,
  input  [63:0] io_in_addr_req_bits_addr,
  input         io_in_addr_req_bits_ce,
  input         io_in_addr_req_bits_we,
  output        io_in_rdata_rep_valid,
  output [63:0] io_in_rdata_rep_bits_rdata,
  input  [63:0] io_in_wdata_req_bits_wdata,
  input  [7:0]  io_in_wdata_req_bits_wmask,
  output        io_in_wdata_rep,
  output        io_out_addr_req_valid,
  output [63:0] io_out_addr_req_bits_addr,
  output        io_out_addr_req_bits_ce,
  output        io_out_addr_req_bits_we,
  input         io_out_rdata_rep_valid,
  input  [63:0] io_out_rdata_rep_bits_rdata,
  output [63:0] io_out_wdata_req_bits_wdata,
  output [7:0]  io_out_wdata_req_bits_wmask,
  input         io_out_wdata_rep
);
  wire  DCACHE_clock; // @[MMIO.scala 12:22]
  wire  DCACHE_reset; // @[MMIO.scala 12:22]
  wire  DCACHE_io_in_addr_req_valid; // @[MMIO.scala 12:22]
  wire [63:0] DCACHE_io_in_addr_req_bits_addr; // @[MMIO.scala 12:22]
  wire  DCACHE_io_in_addr_req_bits_we; // @[MMIO.scala 12:22]
  wire  DCACHE_io_in_rdata_rep_valid; // @[MMIO.scala 12:22]
  wire [63:0] DCACHE_io_in_rdata_rep_bits_rdata; // @[MMIO.scala 12:22]
  wire [63:0] DCACHE_io_in_wdata_req_bits_wdata; // @[MMIO.scala 12:22]
  wire [7:0] DCACHE_io_in_wdata_req_bits_wmask; // @[MMIO.scala 12:22]
  wire  DCACHE_io_in_wdata_rep; // @[MMIO.scala 12:22]
  wire  DCACHE_io_out_addr_req_valid; // @[MMIO.scala 12:22]
  wire [63:0] DCACHE_io_out_addr_req_bits_addr; // @[MMIO.scala 12:22]
  wire  DCACHE_io_out_addr_req_bits_ce; // @[MMIO.scala 12:22]
  wire  DCACHE_io_out_addr_req_bits_we; // @[MMIO.scala 12:22]
  wire  DCACHE_io_out_rdata_rep_valid; // @[MMIO.scala 12:22]
  wire [63:0] DCACHE_io_out_rdata_rep_bits_rdata; // @[MMIO.scala 12:22]
  wire [63:0] DCACHE_io_out_wdata_req_bits_wdata; // @[MMIO.scala 12:22]
  wire  DCACHE_io_out_wdata_rep; // @[MMIO.scala 12:22]
  wire  _GEN_0 = io_in_addr_req_bits_addr >= 64'ha0000000 & io_in_addr_req_bits_addr <= 64'ha2000000 ? 1'h0 :
    io_in_addr_req_valid; // @[MMIO.scala 14:16 19:97 20:35]
  wire  _GEN_1 = io_in_addr_req_bits_addr >= 64'ha0000000 & io_in_addr_req_bits_addr <= 64'ha2000000 ?
    io_in_addr_req_bits_we : DCACHE_io_out_addr_req_bits_we; // @[MMIO.scala 17:10 19:97 22:23]
  wire  _GEN_2 = io_in_addr_req_bits_addr >= 64'ha0000000 & io_in_addr_req_bits_addr <= 64'ha2000000 ?
    io_in_addr_req_bits_ce : DCACHE_io_out_addr_req_bits_ce; // @[MMIO.scala 17:10 19:97 22:23]
  wire [63:0] _GEN_3 = io_in_addr_req_bits_addr >= 64'ha0000000 & io_in_addr_req_bits_addr <= 64'ha2000000 ?
    io_in_addr_req_bits_addr : DCACHE_io_out_addr_req_bits_addr; // @[MMIO.scala 17:10 19:97 22:23]
  wire  _GEN_4 = io_in_addr_req_bits_addr >= 64'ha0000000 & io_in_addr_req_bits_addr <= 64'ha2000000 ?
    io_in_addr_req_valid : DCACHE_io_out_addr_req_valid; // @[MMIO.scala 17:10 19:97 22:23]
  wire  _GEN_6 = io_in_addr_req_bits_addr >= 64'ha0000000 & io_in_addr_req_bits_addr <= 64'ha2000000 ? io_out_wdata_rep
     : DCACHE_io_in_wdata_rep; // @[MMIO.scala 14:16 19:97 23:28]
  wire [63:0] _GEN_7 = io_in_addr_req_bits_addr >= 64'ha0000000 & io_in_addr_req_bits_addr <= 64'ha2000000 ?
    io_out_rdata_rep_bits_rdata : DCACHE_io_in_rdata_rep_bits_rdata; // @[MMIO.scala 14:16 19:97 24:24]
  wire  _GEN_8 = io_in_addr_req_bits_addr >= 64'ha0000000 & io_in_addr_req_bits_addr <= 64'ha2000000 ?
    io_out_rdata_rep_valid : DCACHE_io_in_rdata_rep_valid; // @[MMIO.scala 14:16 19:97 24:24]
  wire [7:0] _GEN_10 = io_in_addr_req_bits_addr >= 64'ha0000000 & io_in_addr_req_bits_addr <= 64'ha2000000 ?
    io_in_wdata_req_bits_wmask : 8'hff; // @[MMIO.scala 17:10 19:97 25:28]
  wire [63:0] _GEN_11 = io_in_addr_req_bits_addr >= 64'ha0000000 & io_in_addr_req_bits_addr <= 64'ha2000000 ?
    io_in_wdata_req_bits_wdata : DCACHE_io_out_wdata_req_bits_wdata; // @[MMIO.scala 17:10 19:97 25:28]
  Cache_1 DCACHE ( // @[MMIO.scala 12:22]
    .clock(DCACHE_clock),
    .reset(DCACHE_reset),
    .io_in_addr_req_valid(DCACHE_io_in_addr_req_valid),
    .io_in_addr_req_bits_addr(DCACHE_io_in_addr_req_bits_addr),
    .io_in_addr_req_bits_we(DCACHE_io_in_addr_req_bits_we),
    .io_in_rdata_rep_valid(DCACHE_io_in_rdata_rep_valid),
    .io_in_rdata_rep_bits_rdata(DCACHE_io_in_rdata_rep_bits_rdata),
    .io_in_wdata_req_bits_wdata(DCACHE_io_in_wdata_req_bits_wdata),
    .io_in_wdata_req_bits_wmask(DCACHE_io_in_wdata_req_bits_wmask),
    .io_in_wdata_rep(DCACHE_io_in_wdata_rep),
    .io_out_addr_req_valid(DCACHE_io_out_addr_req_valid),
    .io_out_addr_req_bits_addr(DCACHE_io_out_addr_req_bits_addr),
    .io_out_addr_req_bits_ce(DCACHE_io_out_addr_req_bits_ce),
    .io_out_addr_req_bits_we(DCACHE_io_out_addr_req_bits_we),
    .io_out_rdata_rep_valid(DCACHE_io_out_rdata_rep_valid),
    .io_out_rdata_rep_bits_rdata(DCACHE_io_out_rdata_rep_bits_rdata),
    .io_out_wdata_req_bits_wdata(DCACHE_io_out_wdata_req_bits_wdata),
    .io_out_wdata_rep(DCACHE_io_out_wdata_rep)
  );
  assign io_in_rdata_rep_valid = io_in_addr_req_valid ? _GEN_8 : DCACHE_io_in_rdata_rep_valid; // @[MMIO.scala 14:16 18:29]
  assign io_in_rdata_rep_bits_rdata = io_in_addr_req_valid ? _GEN_7 : DCACHE_io_in_rdata_rep_bits_rdata; // @[MMIO.scala 14:16 18:29]
  assign io_in_wdata_rep = io_in_addr_req_valid ? _GEN_6 : DCACHE_io_in_wdata_rep; // @[MMIO.scala 14:16 18:29]
  assign io_out_addr_req_valid = io_in_addr_req_valid ? _GEN_4 : DCACHE_io_out_addr_req_valid; // @[MMIO.scala 17:10 18:29]
  assign io_out_addr_req_bits_addr = io_in_addr_req_valid ? _GEN_3 : DCACHE_io_out_addr_req_bits_addr; // @[MMIO.scala 17:10 18:29]
  assign io_out_addr_req_bits_ce = io_in_addr_req_valid ? _GEN_2 : DCACHE_io_out_addr_req_bits_ce; // @[MMIO.scala 17:10 18:29]
  assign io_out_addr_req_bits_we = io_in_addr_req_valid ? _GEN_1 : DCACHE_io_out_addr_req_bits_we; // @[MMIO.scala 17:10 18:29]
  assign io_out_wdata_req_bits_wdata = io_in_addr_req_valid ? _GEN_11 : DCACHE_io_out_wdata_req_bits_wdata; // @[MMIO.scala 17:10 18:29]
  assign io_out_wdata_req_bits_wmask = io_in_addr_req_valid ? _GEN_10 : 8'hff; // @[MMIO.scala 17:10 18:29]
  assign DCACHE_clock = clock;
  assign DCACHE_reset = reset;
  assign DCACHE_io_in_addr_req_valid = io_in_addr_req_valid ? _GEN_0 : io_in_addr_req_valid; // @[MMIO.scala 14:16 18:29]
  assign DCACHE_io_in_addr_req_bits_addr = io_in_addr_req_bits_addr; // @[MMIO.scala 14:16]
  assign DCACHE_io_in_addr_req_bits_we = io_in_addr_req_bits_we; // @[MMIO.scala 14:16]
  assign DCACHE_io_in_wdata_req_bits_wdata = io_in_wdata_req_bits_wdata; // @[MMIO.scala 14:16]
  assign DCACHE_io_in_wdata_req_bits_wmask = io_in_wdata_req_bits_wmask; // @[MMIO.scala 14:16]
  assign DCACHE_io_out_rdata_rep_valid = io_out_rdata_rep_valid; // @[MMIO.scala 17:10]
  assign DCACHE_io_out_rdata_rep_bits_rdata = io_out_rdata_rep_bits_rdata; // @[MMIO.scala 17:10]
  assign DCACHE_io_out_wdata_rep = io_out_wdata_rep; // @[MMIO.scala 17:10]
endmodule
module CoreTop(
  input         clock,
  input         reset,
  output [63:0] io_pc,
  output [31:0] io_inst
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
`endif // RANDOMIZE_REG_INIT
  wire  IF_clock; // @[CoreTop.scala 84:18]
  wire  IF_reset; // @[CoreTop.scala 84:18]
  wire  IF_io_branch_io_is_branch; // @[CoreTop.scala 84:18]
  wire  IF_io_branch_io_is_jump; // @[CoreTop.scala 84:18]
  wire [63:0] IF_io_branch_io_dnpc; // @[CoreTop.scala 84:18]
  wire  IF_io_cache_req_addr_req_valid; // @[CoreTop.scala 84:18]
  wire [63:0] IF_io_cache_req_addr_req_bits_addr; // @[CoreTop.scala 84:18]
  wire  IF_io_cache_req_rdata_rep_ready; // @[CoreTop.scala 84:18]
  wire  IF_io_cache_req_rdata_rep_valid; // @[CoreTop.scala 84:18]
  wire [63:0] IF_io_cache_req_rdata_rep_bits_rdata; // @[CoreTop.scala 84:18]
  wire  IF_io_out_ready; // @[CoreTop.scala 84:18]
  wire  IF_io_out_valid; // @[CoreTop.scala 84:18]
  wire [63:0] IF_io_out_bits_PC; // @[CoreTop.scala 84:18]
  wire [31:0] IF_io_out_bits_Inst; // @[CoreTop.scala 84:18]
  wire  IF_io_flush; // @[CoreTop.scala 84:18]
  wire  ID_io_in_ready; // @[CoreTop.scala 88:18]
  wire  ID_io_in_valid; // @[CoreTop.scala 88:18]
  wire [63:0] ID_io_in_bits_PC; // @[CoreTop.scala 88:18]
  wire [31:0] ID_io_in_bits_Inst; // @[CoreTop.scala 88:18]
  wire [63:0] ID_io_REG1; // @[CoreTop.scala 88:18]
  wire [63:0] ID_io_REG2; // @[CoreTop.scala 88:18]
  wire  ID_io_flush; // @[CoreTop.scala 88:18]
  wire  ID_io_out_ready; // @[CoreTop.scala 88:18]
  wire  ID_io_out_valid; // @[CoreTop.scala 88:18]
  wire [2:0] ID_io_out_bits_ctrl_signal_src1Type; // @[CoreTop.scala 88:18]
  wire [2:0] ID_io_out_bits_ctrl_signal_src2Type; // @[CoreTop.scala 88:18]
  wire [2:0] ID_io_out_bits_ctrl_signal_fuType; // @[CoreTop.scala 88:18]
  wire  ID_io_out_bits_ctrl_signal_inst_valid; // @[CoreTop.scala 88:18]
  wire [4:0] ID_io_out_bits_ctrl_signal_rfSrc1; // @[CoreTop.scala 88:18]
  wire [4:0] ID_io_out_bits_ctrl_signal_rfSrc2; // @[CoreTop.scala 88:18]
  wire  ID_io_out_bits_ctrl_signal_rfWen; // @[CoreTop.scala 88:18]
  wire [6:0] ID_io_out_bits_ctrl_signal_aluoptype; // @[CoreTop.scala 88:18]
  wire [4:0] ID_io_out_bits_ctrl_signal_rfDest; // @[CoreTop.scala 88:18]
  wire [63:0] ID_io_out_bits_ctrl_data_src1; // @[CoreTop.scala 88:18]
  wire [63:0] ID_io_out_bits_ctrl_data_src2; // @[CoreTop.scala 88:18]
  wire [63:0] ID_io_out_bits_ctrl_data_Imm; // @[CoreTop.scala 88:18]
  wire [63:0] ID_io_out_bits_ctrl_flow_PC; // @[CoreTop.scala 88:18]
  wire [31:0] ID_io_out_bits_ctrl_flow_inst; // @[CoreTop.scala 88:18]
  wire  EX_clock; // @[CoreTop.scala 90:18]
  wire  EX_reset; // @[CoreTop.scala 90:18]
  wire  EX_io_in_ready; // @[CoreTop.scala 90:18]
  wire  EX_io_in_valid; // @[CoreTop.scala 90:18]
  wire [2:0] EX_io_in_bits_ctrl_signal_src1Type; // @[CoreTop.scala 90:18]
  wire [2:0] EX_io_in_bits_ctrl_signal_src2Type; // @[CoreTop.scala 90:18]
  wire [2:0] EX_io_in_bits_ctrl_signal_fuType; // @[CoreTop.scala 90:18]
  wire  EX_io_in_bits_ctrl_signal_inst_valid; // @[CoreTop.scala 90:18]
  wire [4:0] EX_io_in_bits_ctrl_signal_rfSrc1; // @[CoreTop.scala 90:18]
  wire [4:0] EX_io_in_bits_ctrl_signal_rfSrc2; // @[CoreTop.scala 90:18]
  wire  EX_io_in_bits_ctrl_signal_rfWen; // @[CoreTop.scala 90:18]
  wire [6:0] EX_io_in_bits_ctrl_signal_aluoptype; // @[CoreTop.scala 90:18]
  wire [4:0] EX_io_in_bits_ctrl_signal_rfDest; // @[CoreTop.scala 90:18]
  wire [63:0] EX_io_in_bits_ctrl_data_src1; // @[CoreTop.scala 90:18]
  wire [63:0] EX_io_in_bits_ctrl_data_src2; // @[CoreTop.scala 90:18]
  wire [63:0] EX_io_in_bits_ctrl_data_Imm; // @[CoreTop.scala 90:18]
  wire [63:0] EX_io_in_bits_ctrl_flow_PC; // @[CoreTop.scala 90:18]
  wire [31:0] EX_io_in_bits_ctrl_flow_inst; // @[CoreTop.scala 90:18]
  wire [63:0] EX_io_src1; // @[CoreTop.scala 90:18]
  wire [63:0] EX_io_src2; // @[CoreTop.scala 90:18]
  wire  EX_io_branchIO_is_branch; // @[CoreTop.scala 90:18]
  wire  EX_io_branchIO_is_jump; // @[CoreTop.scala 90:18]
  wire [63:0] EX_io_branchIO_dnpc; // @[CoreTop.scala 90:18]
  wire  EX_io_out_ready; // @[CoreTop.scala 90:18]
  wire  EX_io_out_valid; // @[CoreTop.scala 90:18]
  wire [2:0] EX_io_out_bits_ctrl_signal_fuType; // @[CoreTop.scala 90:18]
  wire  EX_io_out_bits_ctrl_signal_inst_valid; // @[CoreTop.scala 90:18]
  wire  EX_io_out_bits_ctrl_signal_rfWen; // @[CoreTop.scala 90:18]
  wire [6:0] EX_io_out_bits_ctrl_signal_aluoptype; // @[CoreTop.scala 90:18]
  wire [63:0] EX_io_out_bits_ctrl_flow_PC; // @[CoreTop.scala 90:18]
  wire [31:0] EX_io_out_bits_ctrl_flow_inst; // @[CoreTop.scala 90:18]
  wire [63:0] EX_io_out_bits_ctrl_flow_Dnpc; // @[CoreTop.scala 90:18]
  wire [4:0] EX_io_out_bits_ctrl_rf_rfDest; // @[CoreTop.scala 90:18]
  wire  EX_io_out_bits_ctrl_rf_rfWen; // @[CoreTop.scala 90:18]
  wire [63:0] EX_io_out_bits_ctrl_rf_rfData; // @[CoreTop.scala 90:18]
  wire [63:0] EX_io_out_bits_ctrl_data_src1; // @[CoreTop.scala 90:18]
  wire [63:0] EX_io_out_bits_ctrl_data_src2; // @[CoreTop.scala 90:18]
  wire [63:0] EX_io_out_bits_ctrl_data_Imm; // @[CoreTop.scala 90:18]
  wire  EX_io_is_break; // @[CoreTop.scala 90:18]
  wire  EX_io_is_flush; // @[CoreTop.scala 90:18]
  wire  DIP_is_break; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_0; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_1; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_2; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_3; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_4; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_5; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_6; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_7; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_8; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_9; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_10; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_11; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_12; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_13; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_14; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_15; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_16; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_17; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_18; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_19; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_20; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_21; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_22; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_23; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_24; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_25; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_26; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_27; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_28; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_29; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_30; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_rf_31; // @[CoreTop.scala 92:19]
  wire [31:0] DIP_inst; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_pc; // @[CoreTop.scala 92:19]
  wire  DIP_inst_valid; // @[CoreTop.scala 92:19]
  wire [63:0] DIP_dnpc; // @[CoreTop.scala 92:19]
  wire  DIP_is_skip; // @[CoreTop.scala 92:19]
  reg [63:0] rf [0:31]; // @[RF.scala 7:15]
  wire  rf_bypass_io_Reg1_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_bypass_io_Reg1_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_bypass_io_Reg1_MPORT_data; // @[RF.scala 7:15]
  wire  rf_bypass_io_Reg2_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_bypass_io_Reg2_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_bypass_io_Reg2_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_0_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_0_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_0_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_1_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_1_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_1_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_2_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_2_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_2_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_3_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_3_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_3_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_4_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_4_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_4_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_5_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_5_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_5_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_6_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_6_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_6_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_7_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_7_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_7_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_8_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_8_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_8_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_9_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_9_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_9_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_10_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_10_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_10_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_11_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_11_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_11_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_12_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_12_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_12_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_13_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_13_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_13_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_14_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_14_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_14_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_15_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_15_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_15_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_16_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_16_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_16_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_17_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_17_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_17_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_18_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_18_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_18_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_19_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_19_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_19_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_20_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_20_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_20_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_21_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_21_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_21_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_22_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_22_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_22_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_23_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_23_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_23_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_24_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_24_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_24_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_25_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_25_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_25_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_26_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_26_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_26_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_27_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_27_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_27_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_28_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_28_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_28_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_29_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_29_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_29_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_30_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_30_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_30_MPORT_data; // @[RF.scala 7:15]
  wire  rf_DIP_io_rf_31_MPORT_en; // @[RF.scala 7:15]
  wire [4:0] rf_DIP_io_rf_31_MPORT_addr; // @[RF.scala 7:15]
  wire [63:0] rf_DIP_io_rf_31_MPORT_data; // @[RF.scala 7:15]
  wire [63:0] rf_MPORT_data; // @[RF.scala 7:15]
  wire [4:0] rf_MPORT_addr; // @[RF.scala 7:15]
  wire  rf_MPORT_mask; // @[RF.scala 7:15]
  wire  rf_MPORT_en; // @[RF.scala 7:15]
  wire  MEM_io_in_ready; // @[CoreTop.scala 98:19]
  wire  MEM_io_in_valid; // @[CoreTop.scala 98:19]
  wire [2:0] MEM_io_in_bits_ctrl_signal_fuType; // @[CoreTop.scala 98:19]
  wire  MEM_io_in_bits_ctrl_signal_inst_valid; // @[CoreTop.scala 98:19]
  wire  MEM_io_in_bits_ctrl_signal_rfWen; // @[CoreTop.scala 98:19]
  wire [6:0] MEM_io_in_bits_ctrl_signal_aluoptype; // @[CoreTop.scala 98:19]
  wire [63:0] MEM_io_in_bits_ctrl_flow_PC; // @[CoreTop.scala 98:19]
  wire [31:0] MEM_io_in_bits_ctrl_flow_inst; // @[CoreTop.scala 98:19]
  wire [63:0] MEM_io_in_bits_ctrl_flow_Dnpc; // @[CoreTop.scala 98:19]
  wire [4:0] MEM_io_in_bits_ctrl_rf_rfDest; // @[CoreTop.scala 98:19]
  wire [63:0] MEM_io_in_bits_ctrl_rf_rfData; // @[CoreTop.scala 98:19]
  wire [63:0] MEM_io_in_bits_ctrl_data_src1; // @[CoreTop.scala 98:19]
  wire [63:0] MEM_io_in_bits_ctrl_data_src2; // @[CoreTop.scala 98:19]
  wire [63:0] MEM_io_in_bits_ctrl_data_Imm; // @[CoreTop.scala 98:19]
  wire  MEM_io_out_ready; // @[CoreTop.scala 98:19]
  wire  MEM_io_out_valid; // @[CoreTop.scala 98:19]
  wire  MEM_io_out_bits_ctrl_signal_inst_valid; // @[CoreTop.scala 98:19]
  wire  MEM_io_out_bits_ctrl_signal_rfWen; // @[CoreTop.scala 98:19]
  wire [63:0] MEM_io_out_bits_ctrl_flow_PC; // @[CoreTop.scala 98:19]
  wire [31:0] MEM_io_out_bits_ctrl_flow_inst; // @[CoreTop.scala 98:19]
  wire [63:0] MEM_io_out_bits_ctrl_flow_Dnpc; // @[CoreTop.scala 98:19]
  wire  MEM_io_out_bits_ctrl_flow_skip; // @[CoreTop.scala 98:19]
  wire [4:0] MEM_io_out_bits_ctrl_rf_rfDest; // @[CoreTop.scala 98:19]
  wire  MEM_io_out_bits_ctrl_rf_rfWen; // @[CoreTop.scala 98:19]
  wire [63:0] MEM_io_out_bits_ctrl_rf_rfData; // @[CoreTop.scala 98:19]
  wire  MEM_io_cache_io_addr_req_valid; // @[CoreTop.scala 98:19]
  wire [63:0] MEM_io_cache_io_addr_req_bits_addr; // @[CoreTop.scala 98:19]
  wire  MEM_io_cache_io_addr_req_bits_ce; // @[CoreTop.scala 98:19]
  wire  MEM_io_cache_io_addr_req_bits_we; // @[CoreTop.scala 98:19]
  wire  MEM_io_cache_io_rdata_rep_valid; // @[CoreTop.scala 98:19]
  wire [63:0] MEM_io_cache_io_rdata_rep_bits_rdata; // @[CoreTop.scala 98:19]
  wire [63:0] MEM_io_cache_io_wdata_req_bits_wdata; // @[CoreTop.scala 98:19]
  wire [7:0] MEM_io_cache_io_wdata_req_bits_wmask; // @[CoreTop.scala 98:19]
  wire  MEM_io_cache_io_wdata_rep; // @[CoreTop.scala 98:19]
  wire  WB_io_in_valid; // @[CoreTop.scala 100:18]
  wire  WB_io_in_bits_ctrl_signal_inst_valid; // @[CoreTop.scala 100:18]
  wire  WB_io_in_bits_ctrl_signal_rfWen; // @[CoreTop.scala 100:18]
  wire [63:0] WB_io_in_bits_ctrl_flow_PC; // @[CoreTop.scala 100:18]
  wire [31:0] WB_io_in_bits_ctrl_flow_inst; // @[CoreTop.scala 100:18]
  wire [63:0] WB_io_in_bits_ctrl_flow_Dnpc; // @[CoreTop.scala 100:18]
  wire  WB_io_in_bits_ctrl_flow_skip; // @[CoreTop.scala 100:18]
  wire [4:0] WB_io_in_bits_ctrl_rf_rfDest; // @[CoreTop.scala 100:18]
  wire [63:0] WB_io_in_bits_ctrl_rf_rfData; // @[CoreTop.scala 100:18]
  wire  WB_io_out_ready; // @[CoreTop.scala 100:18]
  wire  WB_io_out_valid; // @[CoreTop.scala 100:18]
  wire  WB_io_out_bits_ctrl_signal_inst_valid; // @[CoreTop.scala 100:18]
  wire [63:0] WB_io_out_bits_ctrl_flow_PC; // @[CoreTop.scala 100:18]
  wire [31:0] WB_io_out_bits_ctrl_flow_inst; // @[CoreTop.scala 100:18]
  wire [63:0] WB_io_out_bits_ctrl_flow_Dnpc; // @[CoreTop.scala 100:18]
  wire  WB_io_out_bits_ctrl_flow_skip; // @[CoreTop.scala 100:18]
  wire [4:0] WB_io_out_bits_ctrl_rf_rfDest; // @[CoreTop.scala 100:18]
  wire  WB_io_out_bits_ctrl_rf_rfWen; // @[CoreTop.scala 100:18]
  wire [63:0] WB_io_out_bits_ctrl_rf_rfData; // @[CoreTop.scala 100:18]
  wire [4:0] bypass_io_EX_rf_rfDest; // @[CoreTop.scala 102:22]
  wire  bypass_io_EX_rf_rfWen; // @[CoreTop.scala 102:22]
  wire [63:0] bypass_io_EX_rf_rfData; // @[CoreTop.scala 102:22]
  wire [4:0] bypass_io_MEM_rf_rfDest; // @[CoreTop.scala 102:22]
  wire  bypass_io_MEM_rf_rfWen; // @[CoreTop.scala 102:22]
  wire [63:0] bypass_io_MEM_rf_rfData; // @[CoreTop.scala 102:22]
  wire [4:0] bypass_io_WB_rf_rfDest; // @[CoreTop.scala 102:22]
  wire  bypass_io_WB_rf_rfWen; // @[CoreTop.scala 102:22]
  wire [63:0] bypass_io_WB_rf_rfData; // @[CoreTop.scala 102:22]
  wire [63:0] bypass_io_Reg1; // @[CoreTop.scala 102:22]
  wire [4:0] bypass_io_reg_index1; // @[CoreTop.scala 102:22]
  wire [63:0] bypass_io_Reg2; // @[CoreTop.scala 102:22]
  wire [4:0] bypass_io_reg_index2; // @[CoreTop.scala 102:22]
  wire [63:0] bypass_io_Bypass_REG1; // @[CoreTop.scala 102:22]
  wire [63:0] bypass_io_Bypass_REG2; // @[CoreTop.scala 102:22]
  wire [4:0] mem_bypass_io_MEM_rf_rfDest; // @[CoreTop.scala 104:25]
  wire  mem_bypass_io_MEM_rf_rfWen; // @[CoreTop.scala 104:25]
  wire [63:0] mem_bypass_io_MEM_rf_rfData; // @[CoreTop.scala 104:25]
  wire [63:0] mem_bypass_io_Reg1; // @[CoreTop.scala 104:25]
  wire [4:0] mem_bypass_io_reg_index1; // @[CoreTop.scala 104:25]
  wire [63:0] mem_bypass_io_Reg2; // @[CoreTop.scala 104:25]
  wire [4:0] mem_bypass_io_reg_index2; // @[CoreTop.scala 104:25]
  wire [63:0] mem_bypass_io_Bypass_REG1; // @[CoreTop.scala 104:25]
  wire [63:0] mem_bypass_io_Bypass_REG2; // @[CoreTop.scala 104:25]
  wire  ICACHE_clock; // @[CoreTop.scala 106:22]
  wire  ICACHE_reset; // @[CoreTop.scala 106:22]
  wire  ICACHE_io_in_addr_req_valid; // @[CoreTop.scala 106:22]
  wire [63:0] ICACHE_io_in_addr_req_bits_addr; // @[CoreTop.scala 106:22]
  wire  ICACHE_io_in_rdata_rep_ready; // @[CoreTop.scala 106:22]
  wire  ICACHE_io_in_rdata_rep_valid; // @[CoreTop.scala 106:22]
  wire [63:0] ICACHE_io_in_rdata_rep_bits_rdata; // @[CoreTop.scala 106:22]
  wire  ICACHE_io_flush; // @[CoreTop.scala 106:22]
  wire  ICACHE_io_out_addr_req_valid; // @[CoreTop.scala 106:22]
  wire [63:0] ICACHE_io_out_addr_req_bits_addr; // @[CoreTop.scala 106:22]
  wire  ICACHE_io_out_addr_req_bits_ce; // @[CoreTop.scala 106:22]
  wire  ICACHE_io_out_rdata_rep_valid; // @[CoreTop.scala 106:22]
  wire [63:0] ICACHE_io_out_rdata_rep_bits_rdata; // @[CoreTop.scala 106:22]
  wire  If_axi_birdge_clock; // @[CoreTop.scala 108:29]
  wire  If_axi_birdge_reset; // @[CoreTop.scala 108:29]
  wire  If_axi_birdge_io_in_addr_req_valid; // @[CoreTop.scala 108:29]
  wire [63:0] If_axi_birdge_io_in_addr_req_bits_addr; // @[CoreTop.scala 108:29]
  wire  If_axi_birdge_io_in_addr_req_bits_ce; // @[CoreTop.scala 108:29]
  wire  If_axi_birdge_io_in_addr_req_bits_we; // @[CoreTop.scala 108:29]
  wire  If_axi_birdge_io_in_rdata_rep_valid; // @[CoreTop.scala 108:29]
  wire [63:0] If_axi_birdge_io_in_rdata_rep_bits_rdata; // @[CoreTop.scala 108:29]
  wire [63:0] If_axi_birdge_io_in_wdata_req_bits_wdata; // @[CoreTop.scala 108:29]
  wire [7:0] If_axi_birdge_io_in_wdata_req_bits_wmask; // @[CoreTop.scala 108:29]
  wire  If_axi_birdge_io_in_wdata_rep; // @[CoreTop.scala 108:29]
  wire  If_axi_birdge_io_out_raddr_req_ready; // @[CoreTop.scala 108:29]
  wire  If_axi_birdge_io_out_raddr_req_valid; // @[CoreTop.scala 108:29]
  wire [63:0] If_axi_birdge_io_out_raddr_req_bits_addr; // @[CoreTop.scala 108:29]
  wire  If_axi_birdge_io_out_waddr_req_ready; // @[CoreTop.scala 108:29]
  wire  If_axi_birdge_io_out_waddr_req_valid; // @[CoreTop.scala 108:29]
  wire [63:0] If_axi_birdge_io_out_waddr_req_bits_addr; // @[CoreTop.scala 108:29]
  wire  If_axi_birdge_io_out_rdata_rep_ready; // @[CoreTop.scala 108:29]
  wire  If_axi_birdge_io_out_rdata_rep_valid; // @[CoreTop.scala 108:29]
  wire [63:0] If_axi_birdge_io_out_rdata_rep_bits_rdata; // @[CoreTop.scala 108:29]
  wire  If_axi_birdge_io_out_wdata_req_valid; // @[CoreTop.scala 108:29]
  wire [63:0] If_axi_birdge_io_out_wdata_req_bits_wdata; // @[CoreTop.scala 108:29]
  wire [7:0] If_axi_birdge_io_out_wdata_req_bits_wmask; // @[CoreTop.scala 108:29]
  wire  If_axi_birdge_io_out_wb_ready; // @[CoreTop.scala 108:29]
  wire  If_axi_birdge_io_out_wb_valid; // @[CoreTop.scala 108:29]
  wire [1:0] If_axi_birdge_io_out_wb_bits; // @[CoreTop.scala 108:29]
  wire  MEM_axi_birdge_clock; // @[CoreTop.scala 109:30]
  wire  MEM_axi_birdge_reset; // @[CoreTop.scala 109:30]
  wire  MEM_axi_birdge_io_in_addr_req_valid; // @[CoreTop.scala 109:30]
  wire [63:0] MEM_axi_birdge_io_in_addr_req_bits_addr; // @[CoreTop.scala 109:30]
  wire  MEM_axi_birdge_io_in_addr_req_bits_ce; // @[CoreTop.scala 109:30]
  wire  MEM_axi_birdge_io_in_addr_req_bits_we; // @[CoreTop.scala 109:30]
  wire  MEM_axi_birdge_io_in_rdata_rep_valid; // @[CoreTop.scala 109:30]
  wire [63:0] MEM_axi_birdge_io_in_rdata_rep_bits_rdata; // @[CoreTop.scala 109:30]
  wire [63:0] MEM_axi_birdge_io_in_wdata_req_bits_wdata; // @[CoreTop.scala 109:30]
  wire [7:0] MEM_axi_birdge_io_in_wdata_req_bits_wmask; // @[CoreTop.scala 109:30]
  wire  MEM_axi_birdge_io_in_wdata_rep; // @[CoreTop.scala 109:30]
  wire  MEM_axi_birdge_io_out_raddr_req_ready; // @[CoreTop.scala 109:30]
  wire  MEM_axi_birdge_io_out_raddr_req_valid; // @[CoreTop.scala 109:30]
  wire [63:0] MEM_axi_birdge_io_out_raddr_req_bits_addr; // @[CoreTop.scala 109:30]
  wire  MEM_axi_birdge_io_out_waddr_req_ready; // @[CoreTop.scala 109:30]
  wire  MEM_axi_birdge_io_out_waddr_req_valid; // @[CoreTop.scala 109:30]
  wire [63:0] MEM_axi_birdge_io_out_waddr_req_bits_addr; // @[CoreTop.scala 109:30]
  wire  MEM_axi_birdge_io_out_rdata_rep_ready; // @[CoreTop.scala 109:30]
  wire  MEM_axi_birdge_io_out_rdata_rep_valid; // @[CoreTop.scala 109:30]
  wire [63:0] MEM_axi_birdge_io_out_rdata_rep_bits_rdata; // @[CoreTop.scala 109:30]
  wire  MEM_axi_birdge_io_out_wdata_req_valid; // @[CoreTop.scala 109:30]
  wire [63:0] MEM_axi_birdge_io_out_wdata_req_bits_wdata; // @[CoreTop.scala 109:30]
  wire [7:0] MEM_axi_birdge_io_out_wdata_req_bits_wmask; // @[CoreTop.scala 109:30]
  wire  MEM_axi_birdge_io_out_wb_ready; // @[CoreTop.scala 109:30]
  wire  MEM_axi_birdge_io_out_wb_valid; // @[CoreTop.scala 109:30]
  wire [1:0] MEM_axi_birdge_io_out_wb_bits; // @[CoreTop.scala 109:30]
  wire  MMEM_reset; // @[CoreTop.scala 112:20]
  wire  MMEM_clk; // @[CoreTop.scala 112:20]
  wire  MMEM_ar_valid; // @[CoreTop.scala 112:20]
  wire  MMEM_ar_ready; // @[CoreTop.scala 112:20]
  wire [63:0] MMEM_araddr; // @[CoreTop.scala 112:20]
  wire  MMEM_r_valid; // @[CoreTop.scala 112:20]
  wire  MMEM_r_ready; // @[CoreTop.scala 112:20]
  wire [63:0] MMEM_rdata; // @[CoreTop.scala 112:20]
  wire  MMEM_aw_valid; // @[CoreTop.scala 112:20]
  wire  MMEM_aw_ready; // @[CoreTop.scala 112:20]
  wire [63:0] MMEM_awaddr; // @[CoreTop.scala 112:20]
  wire  MMEM_w_valid; // @[CoreTop.scala 112:20]
  wire  MMEM_w_ready; // @[CoreTop.scala 112:20]
  wire [63:0] MMEM_wdata; // @[CoreTop.scala 112:20]
  wire [7:0] MMEM_wstrb; // @[CoreTop.scala 112:20]
  wire  MMEM_bvalid; // @[CoreTop.scala 112:20]
  wire  MMEM_bready; // @[CoreTop.scala 112:20]
  wire [1:0] MMEM_bresp; // @[CoreTop.scala 112:20]
  wire  ARBITER_clock; // @[CoreTop.scala 114:23]
  wire  ARBITER_reset; // @[CoreTop.scala 114:23]
  wire  ARBITER_io_in1_raddr_req_ready; // @[CoreTop.scala 114:23]
  wire  ARBITER_io_in1_raddr_req_valid; // @[CoreTop.scala 114:23]
  wire [63:0] ARBITER_io_in1_raddr_req_bits_addr; // @[CoreTop.scala 114:23]
  wire  ARBITER_io_in1_waddr_req_ready; // @[CoreTop.scala 114:23]
  wire  ARBITER_io_in1_waddr_req_valid; // @[CoreTop.scala 114:23]
  wire [63:0] ARBITER_io_in1_waddr_req_bits_addr; // @[CoreTop.scala 114:23]
  wire  ARBITER_io_in1_rdata_rep_valid; // @[CoreTop.scala 114:23]
  wire [63:0] ARBITER_io_in1_rdata_rep_bits_rdata; // @[CoreTop.scala 114:23]
  wire  ARBITER_io_in1_wdata_req_valid; // @[CoreTop.scala 114:23]
  wire [63:0] ARBITER_io_in1_wdata_req_bits_wdata; // @[CoreTop.scala 114:23]
  wire [7:0] ARBITER_io_in1_wdata_req_bits_wmask; // @[CoreTop.scala 114:23]
  wire  ARBITER_io_in1_wb_ready; // @[CoreTop.scala 114:23]
  wire  ARBITER_io_in1_wb_valid; // @[CoreTop.scala 114:23]
  wire [1:0] ARBITER_io_in1_wb_bits; // @[CoreTop.scala 114:23]
  wire  ARBITER_io_in2_raddr_req_ready; // @[CoreTop.scala 114:23]
  wire  ARBITER_io_in2_raddr_req_valid; // @[CoreTop.scala 114:23]
  wire [63:0] ARBITER_io_in2_raddr_req_bits_addr; // @[CoreTop.scala 114:23]
  wire  ARBITER_io_in2_waddr_req_ready; // @[CoreTop.scala 114:23]
  wire  ARBITER_io_in2_waddr_req_valid; // @[CoreTop.scala 114:23]
  wire [63:0] ARBITER_io_in2_waddr_req_bits_addr; // @[CoreTop.scala 114:23]
  wire  ARBITER_io_in2_rdata_rep_valid; // @[CoreTop.scala 114:23]
  wire [63:0] ARBITER_io_in2_rdata_rep_bits_rdata; // @[CoreTop.scala 114:23]
  wire  ARBITER_io_in2_wdata_req_valid; // @[CoreTop.scala 114:23]
  wire [63:0] ARBITER_io_in2_wdata_req_bits_wdata; // @[CoreTop.scala 114:23]
  wire [7:0] ARBITER_io_in2_wdata_req_bits_wmask; // @[CoreTop.scala 114:23]
  wire  ARBITER_io_in2_wb_ready; // @[CoreTop.scala 114:23]
  wire  ARBITER_io_in2_wb_valid; // @[CoreTop.scala 114:23]
  wire [1:0] ARBITER_io_in2_wb_bits; // @[CoreTop.scala 114:23]
  wire  ARBITER_io_out_raddr_req_valid; // @[CoreTop.scala 114:23]
  wire [63:0] ARBITER_io_out_raddr_req_bits_addr; // @[CoreTop.scala 114:23]
  wire  ARBITER_io_out_waddr_req_valid; // @[CoreTop.scala 114:23]
  wire [63:0] ARBITER_io_out_waddr_req_bits_addr; // @[CoreTop.scala 114:23]
  wire  ARBITER_io_out_rdata_rep_valid; // @[CoreTop.scala 114:23]
  wire [63:0] ARBITER_io_out_rdata_rep_bits_rdata; // @[CoreTop.scala 114:23]
  wire  ARBITER_io_out_wdata_req_valid; // @[CoreTop.scala 114:23]
  wire [63:0] ARBITER_io_out_wdata_req_bits_wdata; // @[CoreTop.scala 114:23]
  wire [7:0] ARBITER_io_out_wdata_req_bits_wmask; // @[CoreTop.scala 114:23]
  wire  ARBITER_io_out_wb_ready; // @[CoreTop.scala 114:23]
  wire  ARBITER_io_out_wb_valid; // @[CoreTop.scala 114:23]
  wire [1:0] ARBITER_io_out_wb_bits; // @[CoreTop.scala 114:23]
  wire  MMIO_clock; // @[CoreTop.scala 116:20]
  wire  MMIO_reset; // @[CoreTop.scala 116:20]
  wire  MMIO_io_in_addr_req_valid; // @[CoreTop.scala 116:20]
  wire [63:0] MMIO_io_in_addr_req_bits_addr; // @[CoreTop.scala 116:20]
  wire  MMIO_io_in_addr_req_bits_ce; // @[CoreTop.scala 116:20]
  wire  MMIO_io_in_addr_req_bits_we; // @[CoreTop.scala 116:20]
  wire  MMIO_io_in_rdata_rep_valid; // @[CoreTop.scala 116:20]
  wire [63:0] MMIO_io_in_rdata_rep_bits_rdata; // @[CoreTop.scala 116:20]
  wire [63:0] MMIO_io_in_wdata_req_bits_wdata; // @[CoreTop.scala 116:20]
  wire [7:0] MMIO_io_in_wdata_req_bits_wmask; // @[CoreTop.scala 116:20]
  wire  MMIO_io_in_wdata_rep; // @[CoreTop.scala 116:20]
  wire  MMIO_io_out_addr_req_valid; // @[CoreTop.scala 116:20]
  wire [63:0] MMIO_io_out_addr_req_bits_addr; // @[CoreTop.scala 116:20]
  wire  MMIO_io_out_addr_req_bits_ce; // @[CoreTop.scala 116:20]
  wire  MMIO_io_out_addr_req_bits_we; // @[CoreTop.scala 116:20]
  wire  MMIO_io_out_rdata_rep_valid; // @[CoreTop.scala 116:20]
  wire [63:0] MMIO_io_out_rdata_rep_bits_rdata; // @[CoreTop.scala 116:20]
  wire [63:0] MMIO_io_out_wdata_req_bits_wdata; // @[CoreTop.scala 116:20]
  wire [7:0] MMIO_io_out_wdata_req_bits_wmask; // @[CoreTop.scala 116:20]
  wire  MMIO_io_out_wdata_rep; // @[CoreTop.scala 116:20]
  wire  _T = ID_io_out_ready & ID_io_out_valid; // @[Decoupled.scala 50:35]
  reg  valid; // @[Pipline.scala 8:24]
  wire  _GEN_0 = _T ? 1'h0 : valid; // @[Pipline.scala 10:22 11:13 8:24]
  wire  _T_1 = IF_io_out_valid & ID_io_in_ready; // @[Pipline.scala 13:21]
  wire  _GEN_1 = IF_io_out_valid & ID_io_in_ready | _GEN_0; // @[Pipline.scala 13:37 14:13]
  reg [63:0] ID_io_in_bits_r_PC; // @[Reg.scala 16:16]
  reg [31:0] ID_io_in_bits_r_Inst; // @[Reg.scala 16:16]
  wire  _T_3 = EX_io_out_ready & EX_io_out_valid; // @[Decoupled.scala 50:35]
  reg  valid_1; // @[Pipline.scala 8:24]
  wire  _GEN_5 = _T_3 ? 1'h0 : valid_1; // @[Pipline.scala 10:22 11:13 8:24]
  wire  _T_4 = ID_io_out_valid & EX_io_in_ready; // @[Pipline.scala 13:21]
  wire  _GEN_6 = ID_io_out_valid & EX_io_in_ready | _GEN_5; // @[Pipline.scala 13:37 14:13]
  reg [2:0] EX_io_in_bits_r_ctrl_signal_src1Type; // @[Reg.scala 16:16]
  reg [2:0] EX_io_in_bits_r_ctrl_signal_src2Type; // @[Reg.scala 16:16]
  reg [2:0] EX_io_in_bits_r_ctrl_signal_fuType; // @[Reg.scala 16:16]
  reg  EX_io_in_bits_r_ctrl_signal_inst_valid; // @[Reg.scala 16:16]
  reg [4:0] EX_io_in_bits_r_ctrl_signal_rfSrc1; // @[Reg.scala 16:16]
  reg [4:0] EX_io_in_bits_r_ctrl_signal_rfSrc2; // @[Reg.scala 16:16]
  reg  EX_io_in_bits_r_ctrl_signal_rfWen; // @[Reg.scala 16:16]
  reg [6:0] EX_io_in_bits_r_ctrl_signal_aluoptype; // @[Reg.scala 16:16]
  reg [4:0] EX_io_in_bits_r_ctrl_signal_rfDest; // @[Reg.scala 16:16]
  reg [63:0] EX_io_in_bits_r_ctrl_data_src1; // @[Reg.scala 16:16]
  reg [63:0] EX_io_in_bits_r_ctrl_data_src2; // @[Reg.scala 16:16]
  reg [63:0] EX_io_in_bits_r_ctrl_data_Imm; // @[Reg.scala 16:16]
  reg [63:0] EX_io_in_bits_r_ctrl_flow_PC; // @[Reg.scala 16:16]
  reg [31:0] EX_io_in_bits_r_ctrl_flow_inst; // @[Reg.scala 16:16]
  wire  _T_6 = MEM_io_out_ready & MEM_io_out_valid; // @[Decoupled.scala 50:35]
  reg  valid_2; // @[Pipline.scala 8:24]
  wire  _GEN_24 = _T_6 ? 1'h0 : valid_2; // @[Pipline.scala 10:22 11:13 8:24]
  wire  _T_7 = EX_io_out_valid & MEM_io_in_ready; // @[Pipline.scala 13:21]
  wire  _GEN_25 = EX_io_out_valid & MEM_io_in_ready | _GEN_24; // @[Pipline.scala 13:37 14:13]
  reg [2:0] MEM_io_in_bits_r_ctrl_signal_fuType; // @[Reg.scala 16:16]
  reg  MEM_io_in_bits_r_ctrl_signal_inst_valid; // @[Reg.scala 16:16]
  reg  MEM_io_in_bits_r_ctrl_signal_rfWen; // @[Reg.scala 16:16]
  reg [6:0] MEM_io_in_bits_r_ctrl_signal_aluoptype; // @[Reg.scala 16:16]
  reg [63:0] MEM_io_in_bits_r_ctrl_flow_PC; // @[Reg.scala 16:16]
  reg [31:0] MEM_io_in_bits_r_ctrl_flow_inst; // @[Reg.scala 16:16]
  reg [63:0] MEM_io_in_bits_r_ctrl_flow_Dnpc; // @[Reg.scala 16:16]
  reg [4:0] MEM_io_in_bits_r_ctrl_rf_rfDest; // @[Reg.scala 16:16]
  reg [63:0] MEM_io_in_bits_r_ctrl_rf_rfData; // @[Reg.scala 16:16]
  reg [63:0] MEM_io_in_bits_r_ctrl_data_src1; // @[Reg.scala 16:16]
  reg [63:0] MEM_io_in_bits_r_ctrl_data_src2; // @[Reg.scala 16:16]
  reg [63:0] MEM_io_in_bits_r_ctrl_data_Imm; // @[Reg.scala 16:16]
  wire  _T_9 = WB_io_out_ready & WB_io_out_valid; // @[Decoupled.scala 50:35]
  reg  valid_3; // @[Pipline.scala 8:24]
  wire  _GEN_46 = _T_9 ? 1'h0 : valid_3; // @[Pipline.scala 10:22 11:13 8:24]
  wire  _T_10 = MEM_io_out_valid; // @[Pipline.scala 13:21]
  wire  _GEN_47 = MEM_io_out_valid | _GEN_46; // @[Pipline.scala 13:37 14:13]
  reg  WB_io_in_bits_r_ctrl_signal_inst_valid; // @[Reg.scala 16:16]
  reg  WB_io_in_bits_r_ctrl_signal_rfWen; // @[Reg.scala 16:16]
  reg [63:0] WB_io_in_bits_r_ctrl_flow_PC; // @[Reg.scala 16:16]
  reg [31:0] WB_io_in_bits_r_ctrl_flow_inst; // @[Reg.scala 16:16]
  reg [63:0] WB_io_in_bits_r_ctrl_flow_Dnpc; // @[Reg.scala 16:16]
  reg  WB_io_in_bits_r_ctrl_flow_skip; // @[Reg.scala 16:16]
  reg [4:0] WB_io_in_bits_r_ctrl_rf_rfDest; // @[Reg.scala 16:16]
  reg [63:0] WB_io_in_bits_r_ctrl_rf_rfData; // @[Reg.scala 16:16]
  wire  _T_13 = WB_io_out_bits_ctrl_rf_rfDest == 5'h0; // @[RF.scala 9:61]
  wire [63:0] _T_14 = WB_io_out_bits_ctrl_rf_rfData; // @[RF.scala 9:78]
  reg  DIP_io_is_break_REG; // @[CoreTop.scala 266:37]
  reg  DIP_io_is_break_REG_1; // @[CoreTop.scala 266:29]
  reg [31:0] DIP_io_inst_REG; // @[CoreTop.scala 270:25]
  reg  DIP_io_is_skip_REG; // @[CoreTop.scala 271:28]
  reg  DIP_io_inst_valid_REG; // @[CoreTop.scala 272:31]
  reg [63:0] DIP_io_pc_REG; // @[CoreTop.scala 273:23]
  reg [63:0] DIP_io_dnpc_REG; // @[CoreTop.scala 274:25]
  IF IF ( // @[CoreTop.scala 84:18]
    .clock(IF_clock),
    .reset(IF_reset),
    .io_branch_io_is_branch(IF_io_branch_io_is_branch),
    .io_branch_io_is_jump(IF_io_branch_io_is_jump),
    .io_branch_io_dnpc(IF_io_branch_io_dnpc),
    .io_cache_req_addr_req_valid(IF_io_cache_req_addr_req_valid),
    .io_cache_req_addr_req_bits_addr(IF_io_cache_req_addr_req_bits_addr),
    .io_cache_req_rdata_rep_ready(IF_io_cache_req_rdata_rep_ready),
    .io_cache_req_rdata_rep_valid(IF_io_cache_req_rdata_rep_valid),
    .io_cache_req_rdata_rep_bits_rdata(IF_io_cache_req_rdata_rep_bits_rdata),
    .io_out_ready(IF_io_out_ready),
    .io_out_valid(IF_io_out_valid),
    .io_out_bits_PC(IF_io_out_bits_PC),
    .io_out_bits_Inst(IF_io_out_bits_Inst),
    .io_flush(IF_io_flush)
  );
  ID ID ( // @[CoreTop.scala 88:18]
    .io_in_ready(ID_io_in_ready),
    .io_in_valid(ID_io_in_valid),
    .io_in_bits_PC(ID_io_in_bits_PC),
    .io_in_bits_Inst(ID_io_in_bits_Inst),
    .io_REG1(ID_io_REG1),
    .io_REG2(ID_io_REG2),
    .io_flush(ID_io_flush),
    .io_out_ready(ID_io_out_ready),
    .io_out_valid(ID_io_out_valid),
    .io_out_bits_ctrl_signal_src1Type(ID_io_out_bits_ctrl_signal_src1Type),
    .io_out_bits_ctrl_signal_src2Type(ID_io_out_bits_ctrl_signal_src2Type),
    .io_out_bits_ctrl_signal_fuType(ID_io_out_bits_ctrl_signal_fuType),
    .io_out_bits_ctrl_signal_inst_valid(ID_io_out_bits_ctrl_signal_inst_valid),
    .io_out_bits_ctrl_signal_rfSrc1(ID_io_out_bits_ctrl_signal_rfSrc1),
    .io_out_bits_ctrl_signal_rfSrc2(ID_io_out_bits_ctrl_signal_rfSrc2),
    .io_out_bits_ctrl_signal_rfWen(ID_io_out_bits_ctrl_signal_rfWen),
    .io_out_bits_ctrl_signal_aluoptype(ID_io_out_bits_ctrl_signal_aluoptype),
    .io_out_bits_ctrl_signal_rfDest(ID_io_out_bits_ctrl_signal_rfDest),
    .io_out_bits_ctrl_data_src1(ID_io_out_bits_ctrl_data_src1),
    .io_out_bits_ctrl_data_src2(ID_io_out_bits_ctrl_data_src2),
    .io_out_bits_ctrl_data_Imm(ID_io_out_bits_ctrl_data_Imm),
    .io_out_bits_ctrl_flow_PC(ID_io_out_bits_ctrl_flow_PC),
    .io_out_bits_ctrl_flow_inst(ID_io_out_bits_ctrl_flow_inst)
  );
  EXE EX ( // @[CoreTop.scala 90:18]
    .clock(EX_clock),
    .reset(EX_reset),
    .io_in_ready(EX_io_in_ready),
    .io_in_valid(EX_io_in_valid),
    .io_in_bits_ctrl_signal_src1Type(EX_io_in_bits_ctrl_signal_src1Type),
    .io_in_bits_ctrl_signal_src2Type(EX_io_in_bits_ctrl_signal_src2Type),
    .io_in_bits_ctrl_signal_fuType(EX_io_in_bits_ctrl_signal_fuType),
    .io_in_bits_ctrl_signal_inst_valid(EX_io_in_bits_ctrl_signal_inst_valid),
    .io_in_bits_ctrl_signal_rfSrc1(EX_io_in_bits_ctrl_signal_rfSrc1),
    .io_in_bits_ctrl_signal_rfSrc2(EX_io_in_bits_ctrl_signal_rfSrc2),
    .io_in_bits_ctrl_signal_rfWen(EX_io_in_bits_ctrl_signal_rfWen),
    .io_in_bits_ctrl_signal_aluoptype(EX_io_in_bits_ctrl_signal_aluoptype),
    .io_in_bits_ctrl_signal_rfDest(EX_io_in_bits_ctrl_signal_rfDest),
    .io_in_bits_ctrl_data_src1(EX_io_in_bits_ctrl_data_src1),
    .io_in_bits_ctrl_data_src2(EX_io_in_bits_ctrl_data_src2),
    .io_in_bits_ctrl_data_Imm(EX_io_in_bits_ctrl_data_Imm),
    .io_in_bits_ctrl_flow_PC(EX_io_in_bits_ctrl_flow_PC),
    .io_in_bits_ctrl_flow_inst(EX_io_in_bits_ctrl_flow_inst),
    .io_src1(EX_io_src1),
    .io_src2(EX_io_src2),
    .io_branchIO_is_branch(EX_io_branchIO_is_branch),
    .io_branchIO_is_jump(EX_io_branchIO_is_jump),
    .io_branchIO_dnpc(EX_io_branchIO_dnpc),
    .io_out_ready(EX_io_out_ready),
    .io_out_valid(EX_io_out_valid),
    .io_out_bits_ctrl_signal_fuType(EX_io_out_bits_ctrl_signal_fuType),
    .io_out_bits_ctrl_signal_inst_valid(EX_io_out_bits_ctrl_signal_inst_valid),
    .io_out_bits_ctrl_signal_rfWen(EX_io_out_bits_ctrl_signal_rfWen),
    .io_out_bits_ctrl_signal_aluoptype(EX_io_out_bits_ctrl_signal_aluoptype),
    .io_out_bits_ctrl_flow_PC(EX_io_out_bits_ctrl_flow_PC),
    .io_out_bits_ctrl_flow_inst(EX_io_out_bits_ctrl_flow_inst),
    .io_out_bits_ctrl_flow_Dnpc(EX_io_out_bits_ctrl_flow_Dnpc),
    .io_out_bits_ctrl_rf_rfDest(EX_io_out_bits_ctrl_rf_rfDest),
    .io_out_bits_ctrl_rf_rfWen(EX_io_out_bits_ctrl_rf_rfWen),
    .io_out_bits_ctrl_rf_rfData(EX_io_out_bits_ctrl_rf_rfData),
    .io_out_bits_ctrl_data_src1(EX_io_out_bits_ctrl_data_src1),
    .io_out_bits_ctrl_data_src2(EX_io_out_bits_ctrl_data_src2),
    .io_out_bits_ctrl_data_Imm(EX_io_out_bits_ctrl_data_Imm),
    .io_is_break(EX_io_is_break),
    .io_is_flush(EX_io_is_flush)
  );
  DIP_model DIP ( // @[CoreTop.scala 92:19]
    .is_break(DIP_is_break),
    .rf_0(DIP_rf_0),
    .rf_1(DIP_rf_1),
    .rf_2(DIP_rf_2),
    .rf_3(DIP_rf_3),
    .rf_4(DIP_rf_4),
    .rf_5(DIP_rf_5),
    .rf_6(DIP_rf_6),
    .rf_7(DIP_rf_7),
    .rf_8(DIP_rf_8),
    .rf_9(DIP_rf_9),
    .rf_10(DIP_rf_10),
    .rf_11(DIP_rf_11),
    .rf_12(DIP_rf_12),
    .rf_13(DIP_rf_13),
    .rf_14(DIP_rf_14),
    .rf_15(DIP_rf_15),
    .rf_16(DIP_rf_16),
    .rf_17(DIP_rf_17),
    .rf_18(DIP_rf_18),
    .rf_19(DIP_rf_19),
    .rf_20(DIP_rf_20),
    .rf_21(DIP_rf_21),
    .rf_22(DIP_rf_22),
    .rf_23(DIP_rf_23),
    .rf_24(DIP_rf_24),
    .rf_25(DIP_rf_25),
    .rf_26(DIP_rf_26),
    .rf_27(DIP_rf_27),
    .rf_28(DIP_rf_28),
    .rf_29(DIP_rf_29),
    .rf_30(DIP_rf_30),
    .rf_31(DIP_rf_31),
    .inst(DIP_inst),
    .pc(DIP_pc),
    .inst_valid(DIP_inst_valid),
    .dnpc(DIP_dnpc),
    .is_skip(DIP_is_skip)
  );
  MEM_stage MEM ( // @[CoreTop.scala 98:19]
    .io_in_ready(MEM_io_in_ready),
    .io_in_valid(MEM_io_in_valid),
    .io_in_bits_ctrl_signal_fuType(MEM_io_in_bits_ctrl_signal_fuType),
    .io_in_bits_ctrl_signal_inst_valid(MEM_io_in_bits_ctrl_signal_inst_valid),
    .io_in_bits_ctrl_signal_rfWen(MEM_io_in_bits_ctrl_signal_rfWen),
    .io_in_bits_ctrl_signal_aluoptype(MEM_io_in_bits_ctrl_signal_aluoptype),
    .io_in_bits_ctrl_flow_PC(MEM_io_in_bits_ctrl_flow_PC),
    .io_in_bits_ctrl_flow_inst(MEM_io_in_bits_ctrl_flow_inst),
    .io_in_bits_ctrl_flow_Dnpc(MEM_io_in_bits_ctrl_flow_Dnpc),
    .io_in_bits_ctrl_rf_rfDest(MEM_io_in_bits_ctrl_rf_rfDest),
    .io_in_bits_ctrl_rf_rfData(MEM_io_in_bits_ctrl_rf_rfData),
    .io_in_bits_ctrl_data_src1(MEM_io_in_bits_ctrl_data_src1),
    .io_in_bits_ctrl_data_src2(MEM_io_in_bits_ctrl_data_src2),
    .io_in_bits_ctrl_data_Imm(MEM_io_in_bits_ctrl_data_Imm),
    .io_out_ready(MEM_io_out_ready),
    .io_out_valid(MEM_io_out_valid),
    .io_out_bits_ctrl_signal_inst_valid(MEM_io_out_bits_ctrl_signal_inst_valid),
    .io_out_bits_ctrl_signal_rfWen(MEM_io_out_bits_ctrl_signal_rfWen),
    .io_out_bits_ctrl_flow_PC(MEM_io_out_bits_ctrl_flow_PC),
    .io_out_bits_ctrl_flow_inst(MEM_io_out_bits_ctrl_flow_inst),
    .io_out_bits_ctrl_flow_Dnpc(MEM_io_out_bits_ctrl_flow_Dnpc),
    .io_out_bits_ctrl_flow_skip(MEM_io_out_bits_ctrl_flow_skip),
    .io_out_bits_ctrl_rf_rfDest(MEM_io_out_bits_ctrl_rf_rfDest),
    .io_out_bits_ctrl_rf_rfWen(MEM_io_out_bits_ctrl_rf_rfWen),
    .io_out_bits_ctrl_rf_rfData(MEM_io_out_bits_ctrl_rf_rfData),
    .io_cache_io_addr_req_valid(MEM_io_cache_io_addr_req_valid),
    .io_cache_io_addr_req_bits_addr(MEM_io_cache_io_addr_req_bits_addr),
    .io_cache_io_addr_req_bits_ce(MEM_io_cache_io_addr_req_bits_ce),
    .io_cache_io_addr_req_bits_we(MEM_io_cache_io_addr_req_bits_we),
    .io_cache_io_rdata_rep_valid(MEM_io_cache_io_rdata_rep_valid),
    .io_cache_io_rdata_rep_bits_rdata(MEM_io_cache_io_rdata_rep_bits_rdata),
    .io_cache_io_wdata_req_bits_wdata(MEM_io_cache_io_wdata_req_bits_wdata),
    .io_cache_io_wdata_req_bits_wmask(MEM_io_cache_io_wdata_req_bits_wmask),
    .io_cache_io_wdata_rep(MEM_io_cache_io_wdata_rep)
  );
  WB WB ( // @[CoreTop.scala 100:18]
    .io_in_valid(WB_io_in_valid),
    .io_in_bits_ctrl_signal_inst_valid(WB_io_in_bits_ctrl_signal_inst_valid),
    .io_in_bits_ctrl_signal_rfWen(WB_io_in_bits_ctrl_signal_rfWen),
    .io_in_bits_ctrl_flow_PC(WB_io_in_bits_ctrl_flow_PC),
    .io_in_bits_ctrl_flow_inst(WB_io_in_bits_ctrl_flow_inst),
    .io_in_bits_ctrl_flow_Dnpc(WB_io_in_bits_ctrl_flow_Dnpc),
    .io_in_bits_ctrl_flow_skip(WB_io_in_bits_ctrl_flow_skip),
    .io_in_bits_ctrl_rf_rfDest(WB_io_in_bits_ctrl_rf_rfDest),
    .io_in_bits_ctrl_rf_rfData(WB_io_in_bits_ctrl_rf_rfData),
    .io_out_ready(WB_io_out_ready),
    .io_out_valid(WB_io_out_valid),
    .io_out_bits_ctrl_signal_inst_valid(WB_io_out_bits_ctrl_signal_inst_valid),
    .io_out_bits_ctrl_flow_PC(WB_io_out_bits_ctrl_flow_PC),
    .io_out_bits_ctrl_flow_inst(WB_io_out_bits_ctrl_flow_inst),
    .io_out_bits_ctrl_flow_Dnpc(WB_io_out_bits_ctrl_flow_Dnpc),
    .io_out_bits_ctrl_flow_skip(WB_io_out_bits_ctrl_flow_skip),
    .io_out_bits_ctrl_rf_rfDest(WB_io_out_bits_ctrl_rf_rfDest),
    .io_out_bits_ctrl_rf_rfWen(WB_io_out_bits_ctrl_rf_rfWen),
    .io_out_bits_ctrl_rf_rfData(WB_io_out_bits_ctrl_rf_rfData)
  );
  Bypass bypass ( // @[CoreTop.scala 102:22]
    .io_EX_rf_rfDest(bypass_io_EX_rf_rfDest),
    .io_EX_rf_rfWen(bypass_io_EX_rf_rfWen),
    .io_EX_rf_rfData(bypass_io_EX_rf_rfData),
    .io_MEM_rf_rfDest(bypass_io_MEM_rf_rfDest),
    .io_MEM_rf_rfWen(bypass_io_MEM_rf_rfWen),
    .io_MEM_rf_rfData(bypass_io_MEM_rf_rfData),
    .io_WB_rf_rfDest(bypass_io_WB_rf_rfDest),
    .io_WB_rf_rfWen(bypass_io_WB_rf_rfWen),
    .io_WB_rf_rfData(bypass_io_WB_rf_rfData),
    .io_Reg1(bypass_io_Reg1),
    .io_reg_index1(bypass_io_reg_index1),
    .io_Reg2(bypass_io_Reg2),
    .io_reg_index2(bypass_io_reg_index2),
    .io_Bypass_REG1(bypass_io_Bypass_REG1),
    .io_Bypass_REG2(bypass_io_Bypass_REG2)
  );
  MEM_Bypass mem_bypass ( // @[CoreTop.scala 104:25]
    .io_MEM_rf_rfDest(mem_bypass_io_MEM_rf_rfDest),
    .io_MEM_rf_rfWen(mem_bypass_io_MEM_rf_rfWen),
    .io_MEM_rf_rfData(mem_bypass_io_MEM_rf_rfData),
    .io_Reg1(mem_bypass_io_Reg1),
    .io_reg_index1(mem_bypass_io_reg_index1),
    .io_Reg2(mem_bypass_io_Reg2),
    .io_reg_index2(mem_bypass_io_reg_index2),
    .io_Bypass_REG1(mem_bypass_io_Bypass_REG1),
    .io_Bypass_REG2(mem_bypass_io_Bypass_REG2)
  );
  Cache ICACHE ( // @[CoreTop.scala 106:22]
    .clock(ICACHE_clock),
    .reset(ICACHE_reset),
    .io_in_addr_req_valid(ICACHE_io_in_addr_req_valid),
    .io_in_addr_req_bits_addr(ICACHE_io_in_addr_req_bits_addr),
    .io_in_rdata_rep_ready(ICACHE_io_in_rdata_rep_ready),
    .io_in_rdata_rep_valid(ICACHE_io_in_rdata_rep_valid),
    .io_in_rdata_rep_bits_rdata(ICACHE_io_in_rdata_rep_bits_rdata),
    .io_flush(ICACHE_io_flush),
    .io_out_addr_req_valid(ICACHE_io_out_addr_req_valid),
    .io_out_addr_req_bits_addr(ICACHE_io_out_addr_req_bits_addr),
    .io_out_addr_req_bits_ce(ICACHE_io_out_addr_req_bits_ce),
    .io_out_rdata_rep_valid(ICACHE_io_out_rdata_rep_valid),
    .io_out_rdata_rep_bits_rdata(ICACHE_io_out_rdata_rep_bits_rdata)
  );
  Sram2axi_mulit If_axi_birdge ( // @[CoreTop.scala 108:29]
    .clock(If_axi_birdge_clock),
    .reset(If_axi_birdge_reset),
    .io_in_addr_req_valid(If_axi_birdge_io_in_addr_req_valid),
    .io_in_addr_req_bits_addr(If_axi_birdge_io_in_addr_req_bits_addr),
    .io_in_addr_req_bits_ce(If_axi_birdge_io_in_addr_req_bits_ce),
    .io_in_addr_req_bits_we(If_axi_birdge_io_in_addr_req_bits_we),
    .io_in_rdata_rep_valid(If_axi_birdge_io_in_rdata_rep_valid),
    .io_in_rdata_rep_bits_rdata(If_axi_birdge_io_in_rdata_rep_bits_rdata),
    .io_in_wdata_req_bits_wdata(If_axi_birdge_io_in_wdata_req_bits_wdata),
    .io_in_wdata_req_bits_wmask(If_axi_birdge_io_in_wdata_req_bits_wmask),
    .io_in_wdata_rep(If_axi_birdge_io_in_wdata_rep),
    .io_out_raddr_req_ready(If_axi_birdge_io_out_raddr_req_ready),
    .io_out_raddr_req_valid(If_axi_birdge_io_out_raddr_req_valid),
    .io_out_raddr_req_bits_addr(If_axi_birdge_io_out_raddr_req_bits_addr),
    .io_out_waddr_req_ready(If_axi_birdge_io_out_waddr_req_ready),
    .io_out_waddr_req_valid(If_axi_birdge_io_out_waddr_req_valid),
    .io_out_waddr_req_bits_addr(If_axi_birdge_io_out_waddr_req_bits_addr),
    .io_out_rdata_rep_ready(If_axi_birdge_io_out_rdata_rep_ready),
    .io_out_rdata_rep_valid(If_axi_birdge_io_out_rdata_rep_valid),
    .io_out_rdata_rep_bits_rdata(If_axi_birdge_io_out_rdata_rep_bits_rdata),
    .io_out_wdata_req_valid(If_axi_birdge_io_out_wdata_req_valid),
    .io_out_wdata_req_bits_wdata(If_axi_birdge_io_out_wdata_req_bits_wdata),
    .io_out_wdata_req_bits_wmask(If_axi_birdge_io_out_wdata_req_bits_wmask),
    .io_out_wb_ready(If_axi_birdge_io_out_wb_ready),
    .io_out_wb_valid(If_axi_birdge_io_out_wb_valid),
    .io_out_wb_bits(If_axi_birdge_io_out_wb_bits)
  );
  Sram2axi_mulit MEM_axi_birdge ( // @[CoreTop.scala 109:30]
    .clock(MEM_axi_birdge_clock),
    .reset(MEM_axi_birdge_reset),
    .io_in_addr_req_valid(MEM_axi_birdge_io_in_addr_req_valid),
    .io_in_addr_req_bits_addr(MEM_axi_birdge_io_in_addr_req_bits_addr),
    .io_in_addr_req_bits_ce(MEM_axi_birdge_io_in_addr_req_bits_ce),
    .io_in_addr_req_bits_we(MEM_axi_birdge_io_in_addr_req_bits_we),
    .io_in_rdata_rep_valid(MEM_axi_birdge_io_in_rdata_rep_valid),
    .io_in_rdata_rep_bits_rdata(MEM_axi_birdge_io_in_rdata_rep_bits_rdata),
    .io_in_wdata_req_bits_wdata(MEM_axi_birdge_io_in_wdata_req_bits_wdata),
    .io_in_wdata_req_bits_wmask(MEM_axi_birdge_io_in_wdata_req_bits_wmask),
    .io_in_wdata_rep(MEM_axi_birdge_io_in_wdata_rep),
    .io_out_raddr_req_ready(MEM_axi_birdge_io_out_raddr_req_ready),
    .io_out_raddr_req_valid(MEM_axi_birdge_io_out_raddr_req_valid),
    .io_out_raddr_req_bits_addr(MEM_axi_birdge_io_out_raddr_req_bits_addr),
    .io_out_waddr_req_ready(MEM_axi_birdge_io_out_waddr_req_ready),
    .io_out_waddr_req_valid(MEM_axi_birdge_io_out_waddr_req_valid),
    .io_out_waddr_req_bits_addr(MEM_axi_birdge_io_out_waddr_req_bits_addr),
    .io_out_rdata_rep_ready(MEM_axi_birdge_io_out_rdata_rep_ready),
    .io_out_rdata_rep_valid(MEM_axi_birdge_io_out_rdata_rep_valid),
    .io_out_rdata_rep_bits_rdata(MEM_axi_birdge_io_out_rdata_rep_bits_rdata),
    .io_out_wdata_req_valid(MEM_axi_birdge_io_out_wdata_req_valid),
    .io_out_wdata_req_bits_wdata(MEM_axi_birdge_io_out_wdata_req_bits_wdata),
    .io_out_wdata_req_bits_wmask(MEM_axi_birdge_io_out_wdata_req_bits_wmask),
    .io_out_wb_ready(MEM_axi_birdge_io_out_wb_ready),
    .io_out_wb_valid(MEM_axi_birdge_io_out_wb_valid),
    .io_out_wb_bits(MEM_axi_birdge_io_out_wb_bits)
  );
  SRAM MMEM ( // @[CoreTop.scala 112:20]
    .reset(MMEM_reset),
    .clk(MMEM_clk),
    .ar_valid(MMEM_ar_valid),
    .ar_ready(MMEM_ar_ready),
    .araddr(MMEM_araddr),
    .r_valid(MMEM_r_valid),
    .r_ready(MMEM_r_ready),
    .rdata(MMEM_rdata),
    .aw_valid(MMEM_aw_valid),
    .aw_ready(MMEM_aw_ready),
    .awaddr(MMEM_awaddr),
    .w_valid(MMEM_w_valid),
    .w_ready(MMEM_w_ready),
    .wdata(MMEM_wdata),
    .wstrb(MMEM_wstrb),
    .bvalid(MMEM_bvalid),
    .bready(MMEM_bready),
    .bresp(MMEM_bresp)
  );
  AxiArbiter ARBITER ( // @[CoreTop.scala 114:23]
    .clock(ARBITER_clock),
    .reset(ARBITER_reset),
    .io_in1_raddr_req_ready(ARBITER_io_in1_raddr_req_ready),
    .io_in1_raddr_req_valid(ARBITER_io_in1_raddr_req_valid),
    .io_in1_raddr_req_bits_addr(ARBITER_io_in1_raddr_req_bits_addr),
    .io_in1_waddr_req_ready(ARBITER_io_in1_waddr_req_ready),
    .io_in1_waddr_req_valid(ARBITER_io_in1_waddr_req_valid),
    .io_in1_waddr_req_bits_addr(ARBITER_io_in1_waddr_req_bits_addr),
    .io_in1_rdata_rep_valid(ARBITER_io_in1_rdata_rep_valid),
    .io_in1_rdata_rep_bits_rdata(ARBITER_io_in1_rdata_rep_bits_rdata),
    .io_in1_wdata_req_valid(ARBITER_io_in1_wdata_req_valid),
    .io_in1_wdata_req_bits_wdata(ARBITER_io_in1_wdata_req_bits_wdata),
    .io_in1_wdata_req_bits_wmask(ARBITER_io_in1_wdata_req_bits_wmask),
    .io_in1_wb_ready(ARBITER_io_in1_wb_ready),
    .io_in1_wb_valid(ARBITER_io_in1_wb_valid),
    .io_in1_wb_bits(ARBITER_io_in1_wb_bits),
    .io_in2_raddr_req_ready(ARBITER_io_in2_raddr_req_ready),
    .io_in2_raddr_req_valid(ARBITER_io_in2_raddr_req_valid),
    .io_in2_raddr_req_bits_addr(ARBITER_io_in2_raddr_req_bits_addr),
    .io_in2_waddr_req_ready(ARBITER_io_in2_waddr_req_ready),
    .io_in2_waddr_req_valid(ARBITER_io_in2_waddr_req_valid),
    .io_in2_waddr_req_bits_addr(ARBITER_io_in2_waddr_req_bits_addr),
    .io_in2_rdata_rep_valid(ARBITER_io_in2_rdata_rep_valid),
    .io_in2_rdata_rep_bits_rdata(ARBITER_io_in2_rdata_rep_bits_rdata),
    .io_in2_wdata_req_valid(ARBITER_io_in2_wdata_req_valid),
    .io_in2_wdata_req_bits_wdata(ARBITER_io_in2_wdata_req_bits_wdata),
    .io_in2_wdata_req_bits_wmask(ARBITER_io_in2_wdata_req_bits_wmask),
    .io_in2_wb_ready(ARBITER_io_in2_wb_ready),
    .io_in2_wb_valid(ARBITER_io_in2_wb_valid),
    .io_in2_wb_bits(ARBITER_io_in2_wb_bits),
    .io_out_raddr_req_valid(ARBITER_io_out_raddr_req_valid),
    .io_out_raddr_req_bits_addr(ARBITER_io_out_raddr_req_bits_addr),
    .io_out_waddr_req_valid(ARBITER_io_out_waddr_req_valid),
    .io_out_waddr_req_bits_addr(ARBITER_io_out_waddr_req_bits_addr),
    .io_out_rdata_rep_valid(ARBITER_io_out_rdata_rep_valid),
    .io_out_rdata_rep_bits_rdata(ARBITER_io_out_rdata_rep_bits_rdata),
    .io_out_wdata_req_valid(ARBITER_io_out_wdata_req_valid),
    .io_out_wdata_req_bits_wdata(ARBITER_io_out_wdata_req_bits_wdata),
    .io_out_wdata_req_bits_wmask(ARBITER_io_out_wdata_req_bits_wmask),
    .io_out_wb_ready(ARBITER_io_out_wb_ready),
    .io_out_wb_valid(ARBITER_io_out_wb_valid),
    .io_out_wb_bits(ARBITER_io_out_wb_bits)
  );
  MMIO MMIO ( // @[CoreTop.scala 116:20]
    .clock(MMIO_clock),
    .reset(MMIO_reset),
    .io_in_addr_req_valid(MMIO_io_in_addr_req_valid),
    .io_in_addr_req_bits_addr(MMIO_io_in_addr_req_bits_addr),
    .io_in_addr_req_bits_ce(MMIO_io_in_addr_req_bits_ce),
    .io_in_addr_req_bits_we(MMIO_io_in_addr_req_bits_we),
    .io_in_rdata_rep_valid(MMIO_io_in_rdata_rep_valid),
    .io_in_rdata_rep_bits_rdata(MMIO_io_in_rdata_rep_bits_rdata),
    .io_in_wdata_req_bits_wdata(MMIO_io_in_wdata_req_bits_wdata),
    .io_in_wdata_req_bits_wmask(MMIO_io_in_wdata_req_bits_wmask),
    .io_in_wdata_rep(MMIO_io_in_wdata_rep),
    .io_out_addr_req_valid(MMIO_io_out_addr_req_valid),
    .io_out_addr_req_bits_addr(MMIO_io_out_addr_req_bits_addr),
    .io_out_addr_req_bits_ce(MMIO_io_out_addr_req_bits_ce),
    .io_out_addr_req_bits_we(MMIO_io_out_addr_req_bits_we),
    .io_out_rdata_rep_valid(MMIO_io_out_rdata_rep_valid),
    .io_out_rdata_rep_bits_rdata(MMIO_io_out_rdata_rep_bits_rdata),
    .io_out_wdata_req_bits_wdata(MMIO_io_out_wdata_req_bits_wdata),
    .io_out_wdata_req_bits_wmask(MMIO_io_out_wdata_req_bits_wmask),
    .io_out_wdata_rep(MMIO_io_out_wdata_rep)
  );
  assign rf_bypass_io_Reg1_MPORT_en = 1'h1;
  assign rf_bypass_io_Reg1_MPORT_addr = ID_io_out_bits_ctrl_signal_rfSrc1;
  assign rf_bypass_io_Reg1_MPORT_data = rf[rf_bypass_io_Reg1_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_bypass_io_Reg2_MPORT_en = 1'h1;
  assign rf_bypass_io_Reg2_MPORT_addr = ID_io_out_bits_ctrl_signal_rfSrc2;
  assign rf_bypass_io_Reg2_MPORT_data = rf[rf_bypass_io_Reg2_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_0_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_0_MPORT_addr = 5'h0;
  assign rf_DIP_io_rf_0_MPORT_data = rf[rf_DIP_io_rf_0_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_1_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_1_MPORT_addr = 5'h1;
  assign rf_DIP_io_rf_1_MPORT_data = rf[rf_DIP_io_rf_1_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_2_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_2_MPORT_addr = 5'h2;
  assign rf_DIP_io_rf_2_MPORT_data = rf[rf_DIP_io_rf_2_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_3_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_3_MPORT_addr = 5'h3;
  assign rf_DIP_io_rf_3_MPORT_data = rf[rf_DIP_io_rf_3_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_4_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_4_MPORT_addr = 5'h4;
  assign rf_DIP_io_rf_4_MPORT_data = rf[rf_DIP_io_rf_4_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_5_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_5_MPORT_addr = 5'h5;
  assign rf_DIP_io_rf_5_MPORT_data = rf[rf_DIP_io_rf_5_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_6_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_6_MPORT_addr = 5'h6;
  assign rf_DIP_io_rf_6_MPORT_data = rf[rf_DIP_io_rf_6_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_7_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_7_MPORT_addr = 5'h7;
  assign rf_DIP_io_rf_7_MPORT_data = rf[rf_DIP_io_rf_7_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_8_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_8_MPORT_addr = 5'h8;
  assign rf_DIP_io_rf_8_MPORT_data = rf[rf_DIP_io_rf_8_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_9_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_9_MPORT_addr = 5'h9;
  assign rf_DIP_io_rf_9_MPORT_data = rf[rf_DIP_io_rf_9_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_10_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_10_MPORT_addr = 5'ha;
  assign rf_DIP_io_rf_10_MPORT_data = rf[rf_DIP_io_rf_10_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_11_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_11_MPORT_addr = 5'hb;
  assign rf_DIP_io_rf_11_MPORT_data = rf[rf_DIP_io_rf_11_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_12_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_12_MPORT_addr = 5'hc;
  assign rf_DIP_io_rf_12_MPORT_data = rf[rf_DIP_io_rf_12_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_13_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_13_MPORT_addr = 5'hd;
  assign rf_DIP_io_rf_13_MPORT_data = rf[rf_DIP_io_rf_13_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_14_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_14_MPORT_addr = 5'he;
  assign rf_DIP_io_rf_14_MPORT_data = rf[rf_DIP_io_rf_14_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_15_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_15_MPORT_addr = 5'hf;
  assign rf_DIP_io_rf_15_MPORT_data = rf[rf_DIP_io_rf_15_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_16_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_16_MPORT_addr = 5'h10;
  assign rf_DIP_io_rf_16_MPORT_data = rf[rf_DIP_io_rf_16_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_17_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_17_MPORT_addr = 5'h11;
  assign rf_DIP_io_rf_17_MPORT_data = rf[rf_DIP_io_rf_17_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_18_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_18_MPORT_addr = 5'h12;
  assign rf_DIP_io_rf_18_MPORT_data = rf[rf_DIP_io_rf_18_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_19_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_19_MPORT_addr = 5'h13;
  assign rf_DIP_io_rf_19_MPORT_data = rf[rf_DIP_io_rf_19_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_20_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_20_MPORT_addr = 5'h14;
  assign rf_DIP_io_rf_20_MPORT_data = rf[rf_DIP_io_rf_20_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_21_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_21_MPORT_addr = 5'h15;
  assign rf_DIP_io_rf_21_MPORT_data = rf[rf_DIP_io_rf_21_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_22_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_22_MPORT_addr = 5'h16;
  assign rf_DIP_io_rf_22_MPORT_data = rf[rf_DIP_io_rf_22_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_23_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_23_MPORT_addr = 5'h17;
  assign rf_DIP_io_rf_23_MPORT_data = rf[rf_DIP_io_rf_23_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_24_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_24_MPORT_addr = 5'h18;
  assign rf_DIP_io_rf_24_MPORT_data = rf[rf_DIP_io_rf_24_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_25_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_25_MPORT_addr = 5'h19;
  assign rf_DIP_io_rf_25_MPORT_data = rf[rf_DIP_io_rf_25_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_26_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_26_MPORT_addr = 5'h1a;
  assign rf_DIP_io_rf_26_MPORT_data = rf[rf_DIP_io_rf_26_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_27_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_27_MPORT_addr = 5'h1b;
  assign rf_DIP_io_rf_27_MPORT_data = rf[rf_DIP_io_rf_27_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_28_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_28_MPORT_addr = 5'h1c;
  assign rf_DIP_io_rf_28_MPORT_data = rf[rf_DIP_io_rf_28_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_29_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_29_MPORT_addr = 5'h1d;
  assign rf_DIP_io_rf_29_MPORT_data = rf[rf_DIP_io_rf_29_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_30_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_30_MPORT_addr = 5'h1e;
  assign rf_DIP_io_rf_30_MPORT_data = rf[rf_DIP_io_rf_30_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_DIP_io_rf_31_MPORT_en = 1'h1;
  assign rf_DIP_io_rf_31_MPORT_addr = 5'h1f;
  assign rf_DIP_io_rf_31_MPORT_data = rf[rf_DIP_io_rf_31_MPORT_addr]; // @[RF.scala 7:15]
  assign rf_MPORT_data = _T_13 ? 64'h0 : _T_14;
  assign rf_MPORT_addr = WB_io_out_bits_ctrl_rf_rfDest;
  assign rf_MPORT_mask = 1'h1;
  assign rf_MPORT_en = WB_io_out_bits_ctrl_rf_rfWen;
  assign io_pc = IF_io_out_bits_PC; // @[CoreTop.scala 276:9]
  assign io_inst = WB_io_out_bits_ctrl_flow_inst; // @[CoreTop.scala 275:11]
  assign IF_clock = clock;
  assign IF_reset = reset;
  assign IF_io_branch_io_is_branch = EX_io_branchIO_is_branch; // @[CoreTop.scala 201:19]
  assign IF_io_branch_io_is_jump = EX_io_branchIO_is_jump; // @[CoreTop.scala 201:19]
  assign IF_io_branch_io_dnpc = EX_io_branchIO_dnpc; // @[CoreTop.scala 201:19]
  assign IF_io_cache_req_rdata_rep_valid = ICACHE_io_in_rdata_rep_valid; // @[CoreTop.scala 132:29]
  assign IF_io_cache_req_rdata_rep_bits_rdata = ICACHE_io_in_rdata_rep_bits_rdata; // @[CoreTop.scala 132:29]
  assign IF_io_out_ready = ID_io_in_ready; // @[Pipline.scala 20:16]
  assign IF_io_flush = EX_io_is_flush; // @[CoreTop.scala 189:15]
  assign ID_io_in_valid = valid; // @[Pipline.scala 23:17]
  assign ID_io_in_bits_PC = ID_io_in_bits_r_PC; // @[Pipline.scala 21:16]
  assign ID_io_in_bits_Inst = ID_io_in_bits_r_Inst; // @[Pipline.scala 21:16]
  assign ID_io_REG1 = bypass_io_Bypass_REG1; // @[CoreTop.scala 193:14]
  assign ID_io_REG2 = bypass_io_Bypass_REG2; // @[CoreTop.scala 194:14]
  assign ID_io_flush = EX_io_is_flush; // @[CoreTop.scala 195:15]
  assign ID_io_out_ready = EX_io_in_ready; // @[Pipline.scala 20:16]
  assign EX_clock = clock;
  assign EX_reset = reset;
  assign EX_io_in_valid = valid_1; // @[Pipline.scala 23:17]
  assign EX_io_in_bits_ctrl_signal_src1Type = EX_io_in_bits_r_ctrl_signal_src1Type; // @[Pipline.scala 21:16]
  assign EX_io_in_bits_ctrl_signal_src2Type = EX_io_in_bits_r_ctrl_signal_src2Type; // @[Pipline.scala 21:16]
  assign EX_io_in_bits_ctrl_signal_fuType = EX_io_in_bits_r_ctrl_signal_fuType; // @[Pipline.scala 21:16]
  assign EX_io_in_bits_ctrl_signal_inst_valid = EX_io_in_bits_r_ctrl_signal_inst_valid; // @[Pipline.scala 21:16]
  assign EX_io_in_bits_ctrl_signal_rfSrc1 = EX_io_in_bits_r_ctrl_signal_rfSrc1; // @[Pipline.scala 21:16]
  assign EX_io_in_bits_ctrl_signal_rfSrc2 = EX_io_in_bits_r_ctrl_signal_rfSrc2; // @[Pipline.scala 21:16]
  assign EX_io_in_bits_ctrl_signal_rfWen = EX_io_in_bits_r_ctrl_signal_rfWen; // @[Pipline.scala 21:16]
  assign EX_io_in_bits_ctrl_signal_aluoptype = EX_io_in_bits_r_ctrl_signal_aluoptype; // @[Pipline.scala 21:16]
  assign EX_io_in_bits_ctrl_signal_rfDest = EX_io_in_bits_r_ctrl_signal_rfDest; // @[Pipline.scala 21:16]
  assign EX_io_in_bits_ctrl_data_src1 = EX_io_in_bits_r_ctrl_data_src1; // @[Pipline.scala 21:16]
  assign EX_io_in_bits_ctrl_data_src2 = EX_io_in_bits_r_ctrl_data_src2; // @[Pipline.scala 21:16]
  assign EX_io_in_bits_ctrl_data_Imm = EX_io_in_bits_r_ctrl_data_Imm; // @[Pipline.scala 21:16]
  assign EX_io_in_bits_ctrl_flow_PC = EX_io_in_bits_r_ctrl_flow_PC; // @[Pipline.scala 21:16]
  assign EX_io_in_bits_ctrl_flow_inst = EX_io_in_bits_r_ctrl_flow_inst; // @[Pipline.scala 21:16]
  assign EX_io_src1 = mem_bypass_io_Bypass_REG1; // @[CoreTop.scala 209:14]
  assign EX_io_src2 = mem_bypass_io_Bypass_REG2; // @[CoreTop.scala 210:14]
  assign EX_io_out_ready = MEM_io_in_ready; // @[Pipline.scala 20:16]
  assign DIP_is_break = DIP_io_is_break_REG_1; // @[CoreTop.scala 266:19]
  assign DIP_rf_0 = rf_DIP_io_rf_0_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_1 = rf_DIP_io_rf_1_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_2 = rf_DIP_io_rf_2_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_3 = rf_DIP_io_rf_3_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_4 = rf_DIP_io_rf_4_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_5 = rf_DIP_io_rf_5_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_6 = rf_DIP_io_rf_6_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_7 = rf_DIP_io_rf_7_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_8 = rf_DIP_io_rf_8_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_9 = rf_DIP_io_rf_9_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_10 = rf_DIP_io_rf_10_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_11 = rf_DIP_io_rf_11_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_12 = rf_DIP_io_rf_12_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_13 = rf_DIP_io_rf_13_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_14 = rf_DIP_io_rf_14_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_15 = rf_DIP_io_rf_15_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_16 = rf_DIP_io_rf_16_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_17 = rf_DIP_io_rf_17_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_18 = rf_DIP_io_rf_18_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_19 = rf_DIP_io_rf_19_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_20 = rf_DIP_io_rf_20_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_21 = rf_DIP_io_rf_21_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_22 = rf_DIP_io_rf_22_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_23 = rf_DIP_io_rf_23_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_24 = rf_DIP_io_rf_24_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_25 = rf_DIP_io_rf_25_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_26 = rf_DIP_io_rf_26_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_27 = rf_DIP_io_rf_27_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_28 = rf_DIP_io_rf_28_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_29 = rf_DIP_io_rf_29_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_30 = rf_DIP_io_rf_30_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_rf_31 = rf_DIP_io_rf_31_MPORT_data; // @[CoreTop.scala 268:18]
  assign DIP_inst = DIP_io_inst_REG; // @[CoreTop.scala 270:15]
  assign DIP_pc = DIP_io_pc_REG; // @[CoreTop.scala 273:13]
  assign DIP_inst_valid = DIP_io_inst_valid_REG; // @[CoreTop.scala 272:21]
  assign DIP_dnpc = DIP_io_dnpc_REG; // @[CoreTop.scala 274:15]
  assign DIP_is_skip = DIP_io_is_skip_REG; // @[CoreTop.scala 271:18]
  assign MEM_io_in_valid = valid_2; // @[Pipline.scala 23:17]
  assign MEM_io_in_bits_ctrl_signal_fuType = MEM_io_in_bits_r_ctrl_signal_fuType; // @[Pipline.scala 21:16]
  assign MEM_io_in_bits_ctrl_signal_inst_valid = MEM_io_in_bits_r_ctrl_signal_inst_valid; // @[Pipline.scala 21:16]
  assign MEM_io_in_bits_ctrl_signal_rfWen = MEM_io_in_bits_r_ctrl_signal_rfWen; // @[Pipline.scala 21:16]
  assign MEM_io_in_bits_ctrl_signal_aluoptype = MEM_io_in_bits_r_ctrl_signal_aluoptype; // @[Pipline.scala 21:16]
  assign MEM_io_in_bits_ctrl_flow_PC = MEM_io_in_bits_r_ctrl_flow_PC; // @[Pipline.scala 21:16]
  assign MEM_io_in_bits_ctrl_flow_inst = MEM_io_in_bits_r_ctrl_flow_inst; // @[Pipline.scala 21:16]
  assign MEM_io_in_bits_ctrl_flow_Dnpc = MEM_io_in_bits_r_ctrl_flow_Dnpc; // @[Pipline.scala 21:16]
  assign MEM_io_in_bits_ctrl_rf_rfDest = MEM_io_in_bits_r_ctrl_rf_rfDest; // @[Pipline.scala 21:16]
  assign MEM_io_in_bits_ctrl_rf_rfData = MEM_io_in_bits_r_ctrl_rf_rfData; // @[Pipline.scala 21:16]
  assign MEM_io_in_bits_ctrl_data_src1 = MEM_io_in_bits_r_ctrl_data_src1; // @[Pipline.scala 21:16]
  assign MEM_io_in_bits_ctrl_data_src2 = MEM_io_in_bits_r_ctrl_data_src2; // @[Pipline.scala 21:16]
  assign MEM_io_in_bits_ctrl_data_Imm = MEM_io_in_bits_r_ctrl_data_Imm; // @[Pipline.scala 21:16]
  assign MEM_io_out_ready = 1'h1; // @[Pipline.scala 20:16]
  assign MEM_io_cache_io_rdata_rep_valid = MMIO_io_in_rdata_rep_valid; // @[CoreTop.scala 218:19]
  assign MEM_io_cache_io_rdata_rep_bits_rdata = MMIO_io_in_rdata_rep_bits_rdata; // @[CoreTop.scala 218:19]
  assign MEM_io_cache_io_wdata_rep = MMIO_io_in_wdata_rep; // @[CoreTop.scala 218:19]
  assign WB_io_in_valid = valid_3; // @[Pipline.scala 23:17]
  assign WB_io_in_bits_ctrl_signal_inst_valid = WB_io_in_bits_r_ctrl_signal_inst_valid; // @[Pipline.scala 21:16]
  assign WB_io_in_bits_ctrl_signal_rfWen = WB_io_in_bits_r_ctrl_signal_rfWen; // @[Pipline.scala 21:16]
  assign WB_io_in_bits_ctrl_flow_PC = WB_io_in_bits_r_ctrl_flow_PC; // @[Pipline.scala 21:16]
  assign WB_io_in_bits_ctrl_flow_inst = WB_io_in_bits_r_ctrl_flow_inst; // @[Pipline.scala 21:16]
  assign WB_io_in_bits_ctrl_flow_Dnpc = WB_io_in_bits_r_ctrl_flow_Dnpc; // @[Pipline.scala 21:16]
  assign WB_io_in_bits_ctrl_flow_skip = WB_io_in_bits_r_ctrl_flow_skip; // @[Pipline.scala 21:16]
  assign WB_io_in_bits_ctrl_rf_rfDest = WB_io_in_bits_r_ctrl_rf_rfDest; // @[Pipline.scala 21:16]
  assign WB_io_in_bits_ctrl_rf_rfData = WB_io_in_bits_r_ctrl_rf_rfData; // @[Pipline.scala 21:16]
  assign WB_io_out_ready = 1'h1; // @[CoreTop.scala 262:19]
  assign bypass_io_EX_rf_rfDest = EX_io_out_bits_ctrl_rf_rfDest; // @[CoreTop.scala 202:19]
  assign bypass_io_EX_rf_rfWen = EX_io_out_bits_ctrl_rf_rfWen; // @[CoreTop.scala 202:19]
  assign bypass_io_EX_rf_rfData = EX_io_out_bits_ctrl_rf_rfData; // @[CoreTop.scala 202:19]
  assign bypass_io_MEM_rf_rfDest = MEM_io_out_bits_ctrl_rf_rfDest; // @[CoreTop.scala 252:20]
  assign bypass_io_MEM_rf_rfWen = MEM_io_out_bits_ctrl_rf_rfWen; // @[CoreTop.scala 252:20]
  assign bypass_io_MEM_rf_rfData = MEM_io_out_bits_ctrl_rf_rfData; // @[CoreTop.scala 252:20]
  assign bypass_io_WB_rf_rfDest = WB_io_out_bits_ctrl_rf_rfDest; // @[CoreTop.scala 263:19]
  assign bypass_io_WB_rf_rfWen = WB_io_out_bits_ctrl_rf_rfWen; // @[CoreTop.scala 263:19]
  assign bypass_io_WB_rf_rfData = WB_io_out_bits_ctrl_rf_rfData; // @[CoreTop.scala 263:19]
  assign bypass_io_Reg1 = ID_io_out_bits_ctrl_signal_rfSrc1 == 5'h0 ? 64'h0 : rf_bypass_io_Reg1_MPORT_data; // @[RF.scala 8:37]
  assign bypass_io_reg_index1 = ID_io_out_bits_ctrl_signal_rfSrc1; // @[CoreTop.scala 124:24]
  assign bypass_io_Reg2 = ID_io_out_bits_ctrl_signal_rfSrc2 == 5'h0 ? 64'h0 : rf_bypass_io_Reg2_MPORT_data; // @[RF.scala 8:37]
  assign bypass_io_reg_index2 = ID_io_out_bits_ctrl_signal_rfSrc2; // @[CoreTop.scala 125:24]
  assign mem_bypass_io_MEM_rf_rfDest = MEM_io_out_bits_ctrl_rf_rfDest; // @[CoreTop.scala 254:24]
  assign mem_bypass_io_MEM_rf_rfWen = MEM_io_out_bits_ctrl_rf_rfWen; // @[CoreTop.scala 254:24]
  assign mem_bypass_io_MEM_rf_rfData = MEM_io_out_bits_ctrl_rf_rfData; // @[CoreTop.scala 254:24]
  assign mem_bypass_io_Reg1 = EX_io_in_bits_ctrl_data_src1; // @[CoreTop.scala 204:22]
  assign mem_bypass_io_reg_index1 = EX_io_in_bits_ctrl_signal_rfSrc1; // @[CoreTop.scala 206:28]
  assign mem_bypass_io_Reg2 = EX_io_in_bits_ctrl_data_src2; // @[CoreTop.scala 205:22]
  assign mem_bypass_io_reg_index2 = EX_io_in_bits_ctrl_signal_rfSrc2; // @[CoreTop.scala 207:28]
  assign ICACHE_clock = clock;
  assign ICACHE_reset = reset;
  assign ICACHE_io_in_addr_req_valid = IF_io_cache_req_addr_req_valid; // @[CoreTop.scala 131:28]
  assign ICACHE_io_in_addr_req_bits_addr = IF_io_cache_req_addr_req_bits_addr; // @[CoreTop.scala 131:28]
  assign ICACHE_io_in_rdata_rep_ready = IF_io_cache_req_rdata_rep_ready; // @[CoreTop.scala 132:29]
  assign ICACHE_io_flush = EX_io_is_flush; // @[CoreTop.scala 133:19]
  assign ICACHE_io_out_rdata_rep_valid = If_axi_birdge_io_in_rdata_rep_valid; // @[CoreTop.scala 137:33]
  assign ICACHE_io_out_rdata_rep_bits_rdata = If_axi_birdge_io_in_rdata_rep_bits_rdata; // @[CoreTop.scala 137:33]
  assign If_axi_birdge_clock = clock;
  assign If_axi_birdge_reset = reset;
  assign If_axi_birdge_io_in_addr_req_valid = ICACHE_io_out_addr_req_valid; // @[CoreTop.scala 135:32]
  assign If_axi_birdge_io_in_addr_req_bits_addr = ICACHE_io_out_addr_req_bits_addr; // @[CoreTop.scala 135:32]
  assign If_axi_birdge_io_in_addr_req_bits_ce = ICACHE_io_out_addr_req_bits_ce; // @[CoreTop.scala 135:32]
  assign If_axi_birdge_io_in_addr_req_bits_we = 1'h0; // @[CoreTop.scala 135:32]
  assign If_axi_birdge_io_in_wdata_req_bits_wdata = 64'h0; // @[CoreTop.scala 136:37]
  assign If_axi_birdge_io_in_wdata_req_bits_wmask = 8'h0; // @[CoreTop.scala 136:37]
  assign If_axi_birdge_io_out_raddr_req_ready = ARBITER_io_in2_raddr_req_ready; // @[CoreTop.scala 140:20]
  assign If_axi_birdge_io_out_waddr_req_ready = ARBITER_io_in2_waddr_req_ready; // @[CoreTop.scala 140:20]
  assign If_axi_birdge_io_out_rdata_rep_valid = ARBITER_io_in2_rdata_rep_valid; // @[CoreTop.scala 140:20]
  assign If_axi_birdge_io_out_rdata_rep_bits_rdata = ARBITER_io_in2_rdata_rep_bits_rdata; // @[CoreTop.scala 140:20]
  assign If_axi_birdge_io_out_wb_valid = ARBITER_io_in2_wb_valid; // @[CoreTop.scala 140:20]
  assign If_axi_birdge_io_out_wb_bits = ARBITER_io_in2_wb_bits; // @[CoreTop.scala 140:20]
  assign MEM_axi_birdge_clock = clock;
  assign MEM_axi_birdge_reset = reset;
  assign MEM_axi_birdge_io_in_addr_req_valid = MMIO_io_out_addr_req_valid; // @[CoreTop.scala 224:33]
  assign MEM_axi_birdge_io_in_addr_req_bits_addr = MMIO_io_out_addr_req_bits_addr; // @[CoreTop.scala 224:33]
  assign MEM_axi_birdge_io_in_addr_req_bits_ce = MMIO_io_out_addr_req_bits_ce; // @[CoreTop.scala 224:33]
  assign MEM_axi_birdge_io_in_addr_req_bits_we = MMIO_io_out_addr_req_bits_we; // @[CoreTop.scala 224:33]
  assign MEM_axi_birdge_io_in_wdata_req_bits_wdata = MMIO_io_out_wdata_req_bits_wdata; // @[CoreTop.scala 225:38]
  assign MEM_axi_birdge_io_in_wdata_req_bits_wmask = MMIO_io_out_wdata_req_bits_wmask; // @[CoreTop.scala 225:38]
  assign MEM_axi_birdge_io_out_raddr_req_ready = ARBITER_io_in1_raddr_req_ready; // @[CoreTop.scala 141:20]
  assign MEM_axi_birdge_io_out_waddr_req_ready = ARBITER_io_in1_waddr_req_ready; // @[CoreTop.scala 141:20]
  assign MEM_axi_birdge_io_out_rdata_rep_valid = ARBITER_io_in1_rdata_rep_valid; // @[CoreTop.scala 141:20]
  assign MEM_axi_birdge_io_out_rdata_rep_bits_rdata = ARBITER_io_in1_rdata_rep_bits_rdata; // @[CoreTop.scala 141:20]
  assign MEM_axi_birdge_io_out_wb_valid = ARBITER_io_in1_wb_valid; // @[CoreTop.scala 141:20]
  assign MEM_axi_birdge_io_out_wb_bits = ARBITER_io_in1_wb_bits; // @[CoreTop.scala 141:20]
  assign MMEM_reset = reset; // @[CoreTop.scala 143:19]
  assign MMEM_clk = clock; // @[CoreTop.scala 144:17]
  assign MMEM_ar_valid = ARBITER_io_out_raddr_req_valid; // @[CoreTop.scala 146:22]
  assign MMEM_araddr = ARBITER_io_out_raddr_req_bits_addr; // @[CoreTop.scala 147:20]
  assign MMEM_r_ready = 1'h1; // @[CoreTop.scala 158:21]
  assign MMEM_aw_valid = ARBITER_io_out_waddr_req_valid; // @[CoreTop.scala 150:22]
  assign MMEM_awaddr = ARBITER_io_out_waddr_req_bits_addr; // @[CoreTop.scala 151:20]
  assign MMEM_w_valid = ARBITER_io_out_wdata_req_valid; // @[CoreTop.scala 156:21]
  assign MMEM_wdata = ARBITER_io_out_wdata_req_bits_wdata; // @[CoreTop.scala 154:19]
  assign MMEM_wstrb = ARBITER_io_out_wdata_req_bits_wmask; // @[CoreTop.scala 155:19]
  assign MMEM_bready = ARBITER_io_out_wb_ready; // @[CoreTop.scala 164:20]
  assign ARBITER_clock = clock;
  assign ARBITER_reset = reset;
  assign ARBITER_io_in1_raddr_req_valid = MEM_axi_birdge_io_out_raddr_req_valid; // @[CoreTop.scala 141:20]
  assign ARBITER_io_in1_raddr_req_bits_addr = MEM_axi_birdge_io_out_raddr_req_bits_addr; // @[CoreTop.scala 141:20]
  assign ARBITER_io_in1_waddr_req_valid = MEM_axi_birdge_io_out_waddr_req_valid; // @[CoreTop.scala 141:20]
  assign ARBITER_io_in1_waddr_req_bits_addr = MEM_axi_birdge_io_out_waddr_req_bits_addr; // @[CoreTop.scala 141:20]
  assign ARBITER_io_in1_wdata_req_valid = MEM_axi_birdge_io_out_wdata_req_valid; // @[CoreTop.scala 141:20]
  assign ARBITER_io_in1_wdata_req_bits_wdata = MEM_axi_birdge_io_out_wdata_req_bits_wdata; // @[CoreTop.scala 141:20]
  assign ARBITER_io_in1_wdata_req_bits_wmask = MEM_axi_birdge_io_out_wdata_req_bits_wmask; // @[CoreTop.scala 141:20]
  assign ARBITER_io_in1_wb_ready = MEM_axi_birdge_io_out_wb_ready; // @[CoreTop.scala 141:20]
  assign ARBITER_io_in2_raddr_req_valid = If_axi_birdge_io_out_raddr_req_valid; // @[CoreTop.scala 140:20]
  assign ARBITER_io_in2_raddr_req_bits_addr = If_axi_birdge_io_out_raddr_req_bits_addr; // @[CoreTop.scala 140:20]
  assign ARBITER_io_in2_waddr_req_valid = If_axi_birdge_io_out_waddr_req_valid; // @[CoreTop.scala 140:20]
  assign ARBITER_io_in2_waddr_req_bits_addr = If_axi_birdge_io_out_waddr_req_bits_addr; // @[CoreTop.scala 140:20]
  assign ARBITER_io_in2_wdata_req_valid = If_axi_birdge_io_out_wdata_req_valid; // @[CoreTop.scala 140:20]
  assign ARBITER_io_in2_wdata_req_bits_wdata = If_axi_birdge_io_out_wdata_req_bits_wdata; // @[CoreTop.scala 140:20]
  assign ARBITER_io_in2_wdata_req_bits_wmask = If_axi_birdge_io_out_wdata_req_bits_wmask; // @[CoreTop.scala 140:20]
  assign ARBITER_io_in2_wb_ready = If_axi_birdge_io_out_wb_ready; // @[CoreTop.scala 140:20]
  assign ARBITER_io_out_rdata_rep_valid = MMEM_r_valid; // @[CoreTop.scala 159:36]
  assign ARBITER_io_out_rdata_rep_bits_rdata = MMEM_rdata; // @[CoreTop.scala 160:41]
  assign ARBITER_io_out_wb_valid = MMEM_bvalid; // @[CoreTop.scala 162:29]
  assign ARBITER_io_out_wb_bits = MMEM_bresp; // @[CoreTop.scala 163:28]
  assign MMIO_clock = clock;
  assign MMIO_reset = reset;
  assign MMIO_io_in_addr_req_valid = MEM_io_cache_io_addr_req_valid; // @[CoreTop.scala 218:19]
  assign MMIO_io_in_addr_req_bits_addr = MEM_io_cache_io_addr_req_bits_addr; // @[CoreTop.scala 218:19]
  assign MMIO_io_in_addr_req_bits_ce = MEM_io_cache_io_addr_req_bits_ce; // @[CoreTop.scala 218:19]
  assign MMIO_io_in_addr_req_bits_we = MEM_io_cache_io_addr_req_bits_we; // @[CoreTop.scala 218:19]
  assign MMIO_io_in_wdata_req_bits_wdata = MEM_io_cache_io_wdata_req_bits_wdata; // @[CoreTop.scala 218:19]
  assign MMIO_io_in_wdata_req_bits_wmask = MEM_io_cache_io_wdata_req_bits_wmask; // @[CoreTop.scala 218:19]
  assign MMIO_io_out_rdata_rep_valid = MEM_axi_birdge_io_in_rdata_rep_valid; // @[CoreTop.scala 226:34]
  assign MMIO_io_out_rdata_rep_bits_rdata = MEM_axi_birdge_io_in_rdata_rep_bits_rdata; // @[CoreTop.scala 226:34]
  assign MMIO_io_out_wdata_rep = MEM_axi_birdge_io_in_wdata_rep; // @[CoreTop.scala 227:38]
  always @(posedge clock) begin
    if (rf_MPORT_en & rf_MPORT_mask) begin
      rf[rf_MPORT_addr] <= rf_MPORT_data; // @[RF.scala 7:15]
    end
    if (reset) begin // @[Pipline.scala 8:24]
      valid <= 1'h0; // @[Pipline.scala 8:24]
    end else if (EX_io_is_flush) begin // @[Pipline.scala 16:25]
      valid <= 1'h0; // @[Pipline.scala 17:13]
    end else begin
      valid <= _GEN_1;
    end
    if (_T_1) begin // @[Reg.scala 17:18]
      ID_io_in_bits_r_PC <= IF_io_out_bits_PC; // @[Reg.scala 17:22]
    end
    if (_T_1) begin // @[Reg.scala 17:18]
      ID_io_in_bits_r_Inst <= IF_io_out_bits_Inst; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Pipline.scala 8:24]
      valid_1 <= 1'h0; // @[Pipline.scala 8:24]
    end else if (EX_io_is_flush) begin // @[Pipline.scala 16:25]
      valid_1 <= 1'h0; // @[Pipline.scala 17:13]
    end else begin
      valid_1 <= _GEN_6;
    end
    if (_T_4) begin // @[Reg.scala 17:18]
      EX_io_in_bits_r_ctrl_signal_src1Type <= ID_io_out_bits_ctrl_signal_src1Type; // @[Reg.scala 17:22]
    end
    if (_T_4) begin // @[Reg.scala 17:18]
      EX_io_in_bits_r_ctrl_signal_src2Type <= ID_io_out_bits_ctrl_signal_src2Type; // @[Reg.scala 17:22]
    end
    if (_T_4) begin // @[Reg.scala 17:18]
      EX_io_in_bits_r_ctrl_signal_fuType <= ID_io_out_bits_ctrl_signal_fuType; // @[Reg.scala 17:22]
    end
    if (_T_4) begin // @[Reg.scala 17:18]
      EX_io_in_bits_r_ctrl_signal_inst_valid <= ID_io_out_bits_ctrl_signal_inst_valid; // @[Reg.scala 17:22]
    end
    if (_T_4) begin // @[Reg.scala 17:18]
      EX_io_in_bits_r_ctrl_signal_rfSrc1 <= ID_io_out_bits_ctrl_signal_rfSrc1; // @[Reg.scala 17:22]
    end
    if (_T_4) begin // @[Reg.scala 17:18]
      EX_io_in_bits_r_ctrl_signal_rfSrc2 <= ID_io_out_bits_ctrl_signal_rfSrc2; // @[Reg.scala 17:22]
    end
    if (_T_4) begin // @[Reg.scala 17:18]
      EX_io_in_bits_r_ctrl_signal_rfWen <= ID_io_out_bits_ctrl_signal_rfWen; // @[Reg.scala 17:22]
    end
    if (_T_4) begin // @[Reg.scala 17:18]
      EX_io_in_bits_r_ctrl_signal_aluoptype <= ID_io_out_bits_ctrl_signal_aluoptype; // @[Reg.scala 17:22]
    end
    if (_T_4) begin // @[Reg.scala 17:18]
      EX_io_in_bits_r_ctrl_signal_rfDest <= ID_io_out_bits_ctrl_signal_rfDest; // @[Reg.scala 17:22]
    end
    if (_T_4) begin // @[Reg.scala 17:18]
      EX_io_in_bits_r_ctrl_data_src1 <= ID_io_out_bits_ctrl_data_src1; // @[Reg.scala 17:22]
    end
    if (_T_4) begin // @[Reg.scala 17:18]
      EX_io_in_bits_r_ctrl_data_src2 <= ID_io_out_bits_ctrl_data_src2; // @[Reg.scala 17:22]
    end
    if (_T_4) begin // @[Reg.scala 17:18]
      EX_io_in_bits_r_ctrl_data_Imm <= ID_io_out_bits_ctrl_data_Imm; // @[Reg.scala 17:22]
    end
    if (_T_4) begin // @[Reg.scala 17:18]
      EX_io_in_bits_r_ctrl_flow_PC <= ID_io_out_bits_ctrl_flow_PC; // @[Reg.scala 17:22]
    end
    if (_T_4) begin // @[Reg.scala 17:18]
      EX_io_in_bits_r_ctrl_flow_inst <= ID_io_out_bits_ctrl_flow_inst; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Pipline.scala 8:24]
      valid_2 <= 1'h0; // @[Pipline.scala 8:24]
    end else begin
      valid_2 <= _GEN_25;
    end
    if (_T_7) begin // @[Reg.scala 17:18]
      MEM_io_in_bits_r_ctrl_signal_fuType <= EX_io_out_bits_ctrl_signal_fuType; // @[Reg.scala 17:22]
    end
    if (_T_7) begin // @[Reg.scala 17:18]
      MEM_io_in_bits_r_ctrl_signal_inst_valid <= EX_io_out_bits_ctrl_signal_inst_valid; // @[Reg.scala 17:22]
    end
    if (_T_7) begin // @[Reg.scala 17:18]
      MEM_io_in_bits_r_ctrl_signal_rfWen <= EX_io_out_bits_ctrl_signal_rfWen; // @[Reg.scala 17:22]
    end
    if (_T_7) begin // @[Reg.scala 17:18]
      MEM_io_in_bits_r_ctrl_signal_aluoptype <= EX_io_out_bits_ctrl_signal_aluoptype; // @[Reg.scala 17:22]
    end
    if (_T_7) begin // @[Reg.scala 17:18]
      MEM_io_in_bits_r_ctrl_flow_PC <= EX_io_out_bits_ctrl_flow_PC; // @[Reg.scala 17:22]
    end
    if (_T_7) begin // @[Reg.scala 17:18]
      MEM_io_in_bits_r_ctrl_flow_inst <= EX_io_out_bits_ctrl_flow_inst; // @[Reg.scala 17:22]
    end
    if (_T_7) begin // @[Reg.scala 17:18]
      MEM_io_in_bits_r_ctrl_flow_Dnpc <= EX_io_out_bits_ctrl_flow_Dnpc; // @[Reg.scala 17:22]
    end
    if (_T_7) begin // @[Reg.scala 17:18]
      MEM_io_in_bits_r_ctrl_rf_rfDest <= EX_io_out_bits_ctrl_rf_rfDest; // @[Reg.scala 17:22]
    end
    if (_T_7) begin // @[Reg.scala 17:18]
      MEM_io_in_bits_r_ctrl_rf_rfData <= EX_io_out_bits_ctrl_rf_rfData; // @[Reg.scala 17:22]
    end
    if (_T_7) begin // @[Reg.scala 17:18]
      MEM_io_in_bits_r_ctrl_data_src1 <= EX_io_out_bits_ctrl_data_src1; // @[Reg.scala 17:22]
    end
    if (_T_7) begin // @[Reg.scala 17:18]
      MEM_io_in_bits_r_ctrl_data_src2 <= EX_io_out_bits_ctrl_data_src2; // @[Reg.scala 17:22]
    end
    if (_T_7) begin // @[Reg.scala 17:18]
      MEM_io_in_bits_r_ctrl_data_Imm <= EX_io_out_bits_ctrl_data_Imm; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Pipline.scala 8:24]
      valid_3 <= 1'h0; // @[Pipline.scala 8:24]
    end else begin
      valid_3 <= _GEN_47;
    end
    if (_T_10) begin // @[Reg.scala 17:18]
      WB_io_in_bits_r_ctrl_signal_inst_valid <= MEM_io_out_bits_ctrl_signal_inst_valid; // @[Reg.scala 17:22]
    end
    if (_T_10) begin // @[Reg.scala 17:18]
      WB_io_in_bits_r_ctrl_signal_rfWen <= MEM_io_out_bits_ctrl_signal_rfWen; // @[Reg.scala 17:22]
    end
    if (_T_10) begin // @[Reg.scala 17:18]
      WB_io_in_bits_r_ctrl_flow_PC <= MEM_io_out_bits_ctrl_flow_PC; // @[Reg.scala 17:22]
    end
    if (_T_10) begin // @[Reg.scala 17:18]
      WB_io_in_bits_r_ctrl_flow_inst <= MEM_io_out_bits_ctrl_flow_inst; // @[Reg.scala 17:22]
    end
    if (_T_10) begin // @[Reg.scala 17:18]
      WB_io_in_bits_r_ctrl_flow_Dnpc <= MEM_io_out_bits_ctrl_flow_Dnpc; // @[Reg.scala 17:22]
    end
    if (_T_10) begin // @[Reg.scala 17:18]
      WB_io_in_bits_r_ctrl_flow_skip <= MEM_io_out_bits_ctrl_flow_skip; // @[Reg.scala 17:22]
    end
    if (_T_10) begin // @[Reg.scala 17:18]
      WB_io_in_bits_r_ctrl_rf_rfDest <= MEM_io_out_bits_ctrl_rf_rfDest; // @[Reg.scala 17:22]
    end
    if (_T_10) begin // @[Reg.scala 17:18]
      WB_io_in_bits_r_ctrl_rf_rfData <= MEM_io_out_bits_ctrl_rf_rfData; // @[Reg.scala 17:22]
    end
    DIP_io_is_break_REG <= EX_io_is_break; // @[CoreTop.scala 266:37]
    DIP_io_is_break_REG_1 <= DIP_io_is_break_REG; // @[CoreTop.scala 266:29]
    DIP_io_inst_REG <= WB_io_out_bits_ctrl_flow_inst; // @[CoreTop.scala 270:25]
    DIP_io_is_skip_REG <= WB_io_out_bits_ctrl_flow_skip; // @[CoreTop.scala 271:28]
    DIP_io_inst_valid_REG <= WB_io_out_valid & WB_io_out_bits_ctrl_signal_inst_valid; // @[CoreTop.scala 272:35]
    DIP_io_pc_REG <= WB_io_out_bits_ctrl_flow_PC; // @[CoreTop.scala 273:23]
    DIP_io_dnpc_REG <= WB_io_out_bits_ctrl_flow_Dnpc; // @[CoreTop.scala 274:25]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    rf[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  valid = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  ID_io_in_bits_r_PC = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  ID_io_in_bits_r_Inst = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  valid_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  EX_io_in_bits_r_ctrl_signal_src1Type = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  EX_io_in_bits_r_ctrl_signal_src2Type = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  EX_io_in_bits_r_ctrl_signal_fuType = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  EX_io_in_bits_r_ctrl_signal_inst_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  EX_io_in_bits_r_ctrl_signal_rfSrc1 = _RAND_9[4:0];
  _RAND_10 = {1{`RANDOM}};
  EX_io_in_bits_r_ctrl_signal_rfSrc2 = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  EX_io_in_bits_r_ctrl_signal_rfWen = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  EX_io_in_bits_r_ctrl_signal_aluoptype = _RAND_12[6:0];
  _RAND_13 = {1{`RANDOM}};
  EX_io_in_bits_r_ctrl_signal_rfDest = _RAND_13[4:0];
  _RAND_14 = {2{`RANDOM}};
  EX_io_in_bits_r_ctrl_data_src1 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  EX_io_in_bits_r_ctrl_data_src2 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  EX_io_in_bits_r_ctrl_data_Imm = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  EX_io_in_bits_r_ctrl_flow_PC = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  EX_io_in_bits_r_ctrl_flow_inst = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  valid_2 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  MEM_io_in_bits_r_ctrl_signal_fuType = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  MEM_io_in_bits_r_ctrl_signal_inst_valid = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  MEM_io_in_bits_r_ctrl_signal_rfWen = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  MEM_io_in_bits_r_ctrl_signal_aluoptype = _RAND_23[6:0];
  _RAND_24 = {2{`RANDOM}};
  MEM_io_in_bits_r_ctrl_flow_PC = _RAND_24[63:0];
  _RAND_25 = {1{`RANDOM}};
  MEM_io_in_bits_r_ctrl_flow_inst = _RAND_25[31:0];
  _RAND_26 = {2{`RANDOM}};
  MEM_io_in_bits_r_ctrl_flow_Dnpc = _RAND_26[63:0];
  _RAND_27 = {1{`RANDOM}};
  MEM_io_in_bits_r_ctrl_rf_rfDest = _RAND_27[4:0];
  _RAND_28 = {2{`RANDOM}};
  MEM_io_in_bits_r_ctrl_rf_rfData = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  MEM_io_in_bits_r_ctrl_data_src1 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  MEM_io_in_bits_r_ctrl_data_src2 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  MEM_io_in_bits_r_ctrl_data_Imm = _RAND_31[63:0];
  _RAND_32 = {1{`RANDOM}};
  valid_3 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  WB_io_in_bits_r_ctrl_signal_inst_valid = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  WB_io_in_bits_r_ctrl_signal_rfWen = _RAND_34[0:0];
  _RAND_35 = {2{`RANDOM}};
  WB_io_in_bits_r_ctrl_flow_PC = _RAND_35[63:0];
  _RAND_36 = {1{`RANDOM}};
  WB_io_in_bits_r_ctrl_flow_inst = _RAND_36[31:0];
  _RAND_37 = {2{`RANDOM}};
  WB_io_in_bits_r_ctrl_flow_Dnpc = _RAND_37[63:0];
  _RAND_38 = {1{`RANDOM}};
  WB_io_in_bits_r_ctrl_flow_skip = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  WB_io_in_bits_r_ctrl_rf_rfDest = _RAND_39[4:0];
  _RAND_40 = {2{`RANDOM}};
  WB_io_in_bits_r_ctrl_rf_rfData = _RAND_40[63:0];
  _RAND_41 = {1{`RANDOM}};
  DIP_io_is_break_REG = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  DIP_io_is_break_REG_1 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  DIP_io_inst_REG = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  DIP_io_is_skip_REG = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  DIP_io_inst_valid_REG = _RAND_45[0:0];
  _RAND_46 = {2{`RANDOM}};
  DIP_io_pc_REG = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  DIP_io_dnpc_REG = _RAND_47[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
